-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

entity m2 is
  port (
    clk         : in    std_logic;
    addr        : in    std_logic_vector(10 downto 0);
    data        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of m2 is

  type ROM_ARRAY is array(0 to 2047) of std_logic_vector(7 downto 0);
  constant ROM : ROM_ARRAY := (
    x"C3",x"42",x"F8",x"C3",x"C6",x"F3",x"C3",x"CD", -- 0x0000
    x"F9",x"C3",x"CC",x"F3",x"C3",x"53",x"FA",x"C3", -- 0x0008
    x"34",x"FC",x"C3",x"78",x"FA",x"C3",x"1C",x"F9", -- 0x0010
    x"C3",x"37",x"F9",x"C3",x"EE",x"FA",x"C3",x"63", -- 0x0018
    x"F9",x"C3",x"C9",x"F3",x"C3",x"7F",x"F9",x"C3", -- 0x0020
    x"36",x"F9",x"C3",x"41",x"F9",x"C3",x"EF",x"F8", -- 0x0028
    x"C3",x"6E",x"F9",x"C3",x"6B",x"F9",x"C3",x"78", -- 0x0030
    x"F9",x"C3",x"72",x"F9",x"C3",x"5C",x"F9",x"C3", -- 0x0038
    x"C3",x"F3",x"31",x"C0",x"F3",x"AF",x"D3",x"F8", -- 0x0040
    x"D3",x"F9",x"D3",x"FA",x"32",x"D3",x"F3",x"32", -- 0x0048
    x"D4",x"F3",x"32",x"DE",x"F3",x"3E",x"C3",x"32", -- 0x0050
    x"C6",x"F3",x"32",x"C9",x"F3",x"32",x"CC",x"F3", -- 0x0058
    x"32",x"C3",x"F3",x"21",x"40",x"60",x"22",x"DA", -- 0x0060
    x"F3",x"CD",x"C8",x"F8",x"31",x"C0",x"F3",x"3E", -- 0x0068
    x"8A",x"32",x"03",x"F4",x"3E",x"55",x"32",x"E7", -- 0x0070
    x"F3",x"21",x"6C",x"F8",x"22",x"D8",x"F3",x"AF", -- 0x0078
    x"32",x"E5",x"F3",x"67",x"6F",x"3E",x"90",x"32", -- 0x0080
    x"03",x"F5",x"CD",x"C1",x"F8",x"4F",x"23",x"CD", -- 0x0088
    x"C1",x"F8",x"B9",x"C2",x"AD",x"F8",x"21",x"A6", -- 0x0090
    x"F8",x"CD",x"37",x"F9",x"CD",x"84",x"FA",x"CD", -- 0x0098
    x"7F",x"F9",x"C2",x"96",x"F8",x"E9",x"1F",x"77", -- 0x00A0
    x"77",x"6F",x"64",x"3F",x"00",x"21",x"FF",x"07", -- 0x00A8
    x"11",x"FF",x"BF",x"CD",x"C1",x"F8",x"12",x"1B", -- 0x00B0
    x"2B",x"7C",x"B7",x"F2",x"B3",x"F8",x"C3",x"FD", -- 0x00B8
    x"BF",x"22",x"01",x"F5",x"3A",x"00",x"F5",x"C9", -- 0x00C0
    x"21",x"C0",x"30",x"22",x"CF",x"F3",x"21",x"00", -- 0x00C8
    x"F0",x"22",x"D1",x"F3",x"21",x"37",x"FC",x"22", -- 0x00D0
    x"CD",x"F3",x"22",x"E1",x"F3",x"21",x"36",x"F9", -- 0x00D8
    x"22",x"CA",x"F3",x"21",x"84",x"FA",x"22",x"C7", -- 0x00E0
    x"F3",x"21",x"33",x"FE",x"22",x"C4",x"F3",x"11", -- 0x00E8
    x"4A",x"FE",x"2A",x"D1",x"F3",x"0E",x"07",x"AF", -- 0x00F0
    x"77",x"23",x"1A",x"07",x"07",x"07",x"E6",x"07", -- 0x00F8
    x"47",x"1A",x"E6",x"1F",x"77",x"23",x"0D",x"78", -- 0x0100
    x"A7",x"CA",x"10",x"F9",x"05",x"C3",x"01",x"F9", -- 0x0108
    x"13",x"7A",x"A7",x"C8",x"79",x"A7",x"C2",x"FA", -- 0x0110
    x"F8",x"C3",x"F5",x"F8",x"F5",x"0F",x"0F",x"0F", -- 0x0118
    x"0F",x"CD",x"25",x"F9",x"F1",x"E6",x"0F",x"FE", -- 0x0120
    x"0A",x"FA",x"2E",x"F9",x"C6",x"07",x"C6",x"30", -- 0x0128
    x"C5",x"4F",x"CD",x"09",x"F8",x"C1",x"C9",x"7E", -- 0x0130
    x"A7",x"C8",x"CD",x"30",x"F9",x"23",x"C3",x"37", -- 0x0138
    x"F9",x"01",x"00",x"00",x"79",x"86",x"4F",x"F5", -- 0x0140
    x"CD",x"56",x"F9",x"CA",x"76",x"FA",x"F1",x"78", -- 0x0148
    x"8E",x"47",x"23",x"C3",x"44",x"F9",x"7C",x"BA", -- 0x0150
    x"C0",x"7D",x"BB",x"C9",x"7D",x"07",x"07",x"6F", -- 0x0158
    x"22",x"D6",x"F3",x"2A",x"D6",x"F3",x"7D",x"0F", -- 0x0160
    x"0F",x"6F",x"C9",x"22",x"E3",x"F3",x"2A",x"E3", -- 0x0168
    x"F3",x"C9",x"D3",x"F9",x"71",x"C3",x"7B",x"F9", -- 0x0170
    x"D3",x"F9",x"4E",x"AF",x"D3",x"F9",x"C9",x"3E", -- 0x0178
    x"FF",x"CD",x"B4",x"F9",x"22",x"EE",x"F3",x"EB", -- 0x0180
    x"CD",x"B2",x"F9",x"EB",x"E5",x"CD",x"CB",x"F9", -- 0x0188
    x"77",x"CD",x"56",x"F9",x"23",x"C2",x"8D",x"F9", -- 0x0190
    x"CD",x"CB",x"F9",x"CD",x"B2",x"F9",x"CD",x"B2", -- 0x0198
    x"F9",x"44",x"4D",x"E1",x"C5",x"CD",x"41",x"F9", -- 0x01A0
    x"D1",x"60",x"69",x"CD",x"56",x"F9",x"2A",x"EE", -- 0x01A8
    x"F3",x"C9",x"3E",x"08",x"CD",x"CD",x"F9",x"67", -- 0x01B0
    x"CD",x"CB",x"F9",x"6F",x"C9",x"3A",x"DA",x"F3", -- 0x01B8
    x"C3",x"C6",x"F9",x"3A",x"DB",x"F3",x"3D",x"C2", -- 0x01C0
    x"C6",x"F9",x"C9",x"3E",x"08",x"C5",x"D5",x"E5", -- 0x01C8
    x"0E",x"00",x"57",x"CD",x"45",x"FA",x"5F",x"00", -- 0x01D0
    x"00",x"00",x"00",x"79",x"E6",x"7F",x"07",x"4F", -- 0x01D8
    x"00",x"06",x"00",x"05",x"C2",x"F3",x"F9",x"00", -- 0x01E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01E8
    x"C3",x"4F",x"FA",x"CD",x"45",x"FA",x"BB",x"CA", -- 0x01F0
    x"E3",x"F9",x"00",x"B1",x"4F",x"CD",x"C3",x"F9", -- 0x01F8
    x"CD",x"45",x"FA",x"5F",x"B2",x"F2",x"39",x"FA", -- 0x0200
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0208
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0210
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0218
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3E", -- 0x0220
    x"E6",x"91",x"CA",x"34",x"FA",x"3E",x"19",x"91", -- 0x0228
    x"C2",x"DB",x"F9",x"2F",x"32",x"DC",x"F3",x"16", -- 0x0230
    x"09",x"15",x"C2",x"DB",x"F9",x"3A",x"DC",x"F3", -- 0x0238
    x"A9",x"E1",x"D1",x"C1",x"C9",x"3A",x"02",x"F4", -- 0x0240
    x"0F",x"0F",x"0F",x"0F",x"E6",x"01",x"C9",x"2A", -- 0x0248
    x"D8",x"F3",x"E9",x"F5",x"C5",x"06",x"08",x"00", -- 0x0250
    x"00",x"00",x"00",x"00",x"79",x"07",x"4F",x"3E", -- 0x0258
    x"01",x"A9",x"32",x"02",x"F4",x"CD",x"BD",x"F9", -- 0x0260
    x"3E",x"00",x"A9",x"32",x"02",x"F4",x"CD",x"BD", -- 0x0268
    x"F9",x"05",x"C2",x"5C",x"FA",x"C1",x"F1",x"C9", -- 0x0270
    x"AF",x"32",x"00",x"F4",x"3A",x"01",x"F4",x"3C", -- 0x0278
    x"C8",x"3E",x"FF",x"C9",x"C5",x"D5",x"E5",x"CD", -- 0x0280
    x"EE",x"FA",x"FE",x"FF",x"C2",x"92",x"FA",x"32", -- 0x0288
    x"E6",x"F3",x"16",x"00",x"13",x"1D",x"1C",x"CC", -- 0x0290
    x"72",x"FD",x"CD",x"EE",x"FA",x"3C",x"CA",x"94", -- 0x0298
    x"FA",x"F5",x"7A",x"0F",x"D4",x"72",x"FD",x"F1", -- 0x02A0
    x"3D",x"F2",x"CE",x"FA",x"11",x"40",x"55",x"21", -- 0x02A8
    x"E5",x"F3",x"7E",x"2F",x"77",x"32",x"02",x"F4", -- 0x02B0
    x"A7",x"7A",x"CA",x"BE",x"FA",x"7B",x"32",x"E7", -- 0x02B8
    x"F3",x"CD",x"EE",x"FA",x"3C",x"C2",x"C1",x"FA", -- 0x02C0
    x"CD",x"72",x"FD",x"C3",x"92",x"FA",x"5F",x"16", -- 0x02C8
    x"14",x"21",x"E6",x"F3",x"BE",x"CA",x"E3",x"FA", -- 0x02D0
    x"15",x"CA",x"E3",x"FA",x"CD",x"EE",x"FA",x"BB", -- 0x02D8
    x"CA",x"D8",x"FA",x"CD",x"3F",x"F8",x"73",x"CD", -- 0x02E0
    x"72",x"FD",x"7B",x"C3",x"00",x"FD",x"C5",x"D5", -- 0x02E8
    x"E5",x"21",x"00",x"FD",x"E5",x"06",x"00",x"16", -- 0x02F0
    x"09",x"0E",x"FE",x"79",x"32",x"00",x"F4",x"07", -- 0x02F8
    x"4F",x"3A",x"01",x"F4",x"FE",x"FF",x"CA",x"1A", -- 0x0300
    x"FB",x"5F",x"21",x"00",x"06",x"2B",x"7C",x"B5", -- 0x0308
    x"C2",x"0D",x"FB",x"3A",x"01",x"F4",x"BB",x"CA", -- 0x0310
    x"2D",x"FB",x"78",x"C6",x"08",x"47",x"15",x"C2", -- 0x0318
    x"FB",x"FA",x"3A",x"02",x"F4",x"E6",x"80",x"3E", -- 0x0320
    x"FE",x"C8",x"3C",x"C9",x"04",x"1F",x"DA",x"2C", -- 0x0328
    x"FB",x"78",x"E6",x"3F",x"FE",x"10",x"DA",x"97", -- 0x0330
    x"FB",x"FE",x"3F",x"47",x"3E",x"20",x"C8",x"3A", -- 0x0338
    x"02",x"F4",x"4F",x"E6",x"40",x"C2",x"4C",x"FB", -- 0x0340
    x"78",x"E6",x"1F",x"C9",x"3A",x"E5",x"F3",x"A7", -- 0x0348
    x"C2",x"7B",x"FB",x"79",x"E6",x"20",x"78",x"CA", -- 0x0350
    x"67",x"FB",x"FE",x"1C",x"FA",x"73",x"FB",x"FE", -- 0x0358
    x"20",x"FA",x"75",x"FB",x"C3",x"73",x"FB",x"FE", -- 0x0360
    x"1C",x"DA",x"75",x"FB",x"FE",x"20",x"DA",x"73", -- 0x0368
    x"FB",x"C6",x"20",x"C6",x"10",x"C6",x"10",x"E1", -- 0x0370
    x"C3",x"00",x"FD",x"79",x"E6",x"20",x"78",x"CA", -- 0x0378
    x"8F",x"FB",x"FE",x"1C",x"FA",x"73",x"FB",x"FE", -- 0x0380
    x"20",x"FA",x"75",x"FB",x"C3",x"71",x"FB",x"FE", -- 0x0388
    x"1C",x"FA",x"75",x"FB",x"C3",x"73",x"FB",x"21", -- 0x0390
    x"A0",x"FB",x"4F",x"06",x"00",x"09",x"7E",x"C9", -- 0x0398
    x"0C",x"1F",x"1B",x"00",x"01",x"02",x"03",x"04", -- 0x03A0
    x"09",x"0A",x"0D",x"7F",x"08",x"19",x"18",x"1A", -- 0x03A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"00", -- 0x03B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80", -- 0x03E0
    x"00",x"80",x"00",x"00",x"00",x"00",x"00",x"80", -- 0x03E8
    x"00",x"40",x"00",x"40",x"00",x"00",x"00",x"00", -- 0x03F0
    x"00",x"00",x"00",x"40",x"00",x"40",x"00",x"00", -- 0x03F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0400
    x"00",x"00",x"00",x"40",x"00",x"00",x"00",x"00", -- 0x0408
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0410
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0418
    x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"00", -- 0x0420
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0428
    x"00",x"00",x"00",x"00",x"C5",x"4F",x"06",x"C5", -- 0x0430
    x"D5",x"E5",x"F5",x"79",x"FE",x"1B",x"3E",x"F0", -- 0x0438
    x"CA",x"8A",x"FD",x"3A",x"DE",x"F3",x"A7",x"C2", -- 0x0440
    x"90",x"FD",x"79",x"FE",x"7F",x"C2",x"5A",x"FC", -- 0x0448
    x"3A",x"D3",x"F3",x"2F",x"32",x"D3",x"F3",x"C3", -- 0x0450
    x"FF",x"FC",x"26",x"20",x"94",x"DA",x"A4",x"FC", -- 0x0458
    x"6F",x"29",x"29",x"29",x"EB",x"2A",x"D1",x"F3", -- 0x0460
    x"19",x"EB",x"CD",x"44",x"FD",x"EB",x"3E",x"16", -- 0x0468
    x"F5",x"E5",x"3A",x"D3",x"F3",x"AE",x"E6",x"3F", -- 0x0470
    x"6F",x"3A",x"DD",x"F3",x"3D",x"26",x"00",x"29", -- 0x0478
    x"29",x"3C",x"C2",x"7F",x"FC",x"EB",x"78",x"AE", -- 0x0480
    x"A6",x"B2",x"77",x"24",x"79",x"AE",x"A6",x"B3", -- 0x0488
    x"77",x"25",x"2C",x"EB",x"E1",x"23",x"F1",x"D6", -- 0x0490
    x"03",x"F2",x"70",x"FC",x"21",x"05",x"FD",x"FE", -- 0x0498
    x"F8",x"C2",x"70",x"FC",x"2A",x"D6",x"F3",x"CD", -- 0x04A0
    x"04",x"FD",x"09",x"7C",x"FE",x"19",x"DA",x"FC", -- 0x04A8
    x"FC",x"C2",x"FA",x"FC",x"14",x"62",x"CA",x"FC", -- 0x04B0
    x"FC",x"E5",x"21",x"00",x"00",x"39",x"22",x"DF", -- 0x04B8
    x"F3",x"3A",x"D0",x"F3",x"47",x"3A",x"CF",x"F3", -- 0x04C0
    x"67",x"3A",x"D4",x"F3",x"6F",x"CD",x"6A",x"FD", -- 0x04C8
    x"4F",x"79",x"C6",x"0A",x"6F",x"F9",x"69",x"3E", -- 0x04D0
    x"F0",x"D1",x"73",x"2C",x"72",x"2C",x"D1",x"73", -- 0x04D8
    x"2C",x"72",x"2C",x"BD",x"D2",x"D9",x"FC",x"3A", -- 0x04E0
    x"D3",x"F3",x"33",x"77",x"2C",x"C2",x"EA",x"FC", -- 0x04E8
    x"24",x"05",x"C2",x"D1",x"FC",x"2A",x"DF",x"F3", -- 0x04F0
    x"F9",x"E1",x"26",x"18",x"22",x"D6",x"F3",x"F1", -- 0x04F8
    x"E1",x"D1",x"C1",x"C9",x"01",x"00",x"01",x"51", -- 0x0500
    x"3C",x"CC",x"EC",x"FD",x"CA",x"3F",x"FD",x"FE", -- 0x0508
    x"EB",x"C8",x"15",x"C6",x"05",x"C8",x"14",x"06", -- 0x0510
    x"FF",x"3C",x"C8",x"0E",x"FC",x"FE",x"EF",x"C8", -- 0x0518
    x"01",x"00",x"00",x"FE",x"F0",x"C2",x"2F",x"FD", -- 0x0520
    x"7D",x"E6",x"E0",x"C6",x"20",x"6F",x"C9",x"0E", -- 0x0528
    x"04",x"3C",x"C8",x"FE",x"EF",x"CA",x"3F",x"F8", -- 0x0530
    x"C6",x"0B",x"CA",x"40",x"FD",x"3C",x"C0",x"62", -- 0x0538
    x"6A",x"42",x"4A",x"C9",x"2A",x"D6",x"F3",x"7D", -- 0x0540
    x"0F",x"6F",x"0F",x"85",x"47",x"6C",x"3A",x"CF", -- 0x0548
    x"F3",x"67",x"78",x"25",x"24",x"D6",x"04",x"D2", -- 0x0550
    x"54",x"FD",x"32",x"DD",x"F3",x"E5",x"21",x"FC", -- 0x0558
    x"00",x"29",x"29",x"3C",x"C2",x"61",x"FD",x"44", -- 0x0560
    x"4D",x"E1",x"7D",x"07",x"07",x"07",x"85",x"85", -- 0x0568
    x"6F",x"C9",x"CD",x"44",x"FD",x"C6",x"09",x"6F", -- 0x0570
    x"78",x"AE",x"77",x"24",x"79",x"AE",x"77",x"25", -- 0x0578
    x"C9",x"79",x"FE",x"59",x"C2",x"9E",x"FD",x"3E", -- 0x0580
    x"02",x"B0",x"32",x"DE",x"F3",x"C3",x"FF",x"FC", -- 0x0588
    x"47",x"E6",x"03",x"CA",x"81",x"FD",x"3D",x"CA", -- 0x0590
    x"D3",x"FD",x"3D",x"CA",x"E1",x"FD",x"AF",x"32", -- 0x0598
    x"DE",x"F3",x"79",x"FE",x"4A",x"CA",x"F6",x"FD", -- 0x05A0
    x"FE",x"4B",x"CA",x"1E",x"FE",x"21",x"4A",x"FC", -- 0x05A8
    x"E5",x"0E",x"18",x"FE",x"43",x"C8",x"0C",x"FE", -- 0x05B0
    x"41",x"C8",x"0C",x"FE",x"42",x"C8",x"0E",x"08", -- 0x05B8
    x"FE",x"44",x"C8",x"0E",x"0C",x"FE",x"48",x"C8", -- 0x05C0
    x"0E",x"1F",x"FE",x"45",x"C8",x"B9",x"C8",x"E1", -- 0x05C8
    x"C3",x"FF",x"FC",x"79",x"D6",x"20",x"07",x"07", -- 0x05D0
    x"E6",x"FC",x"32",x"D6",x"F3",x"AF",x"C3",x"8A", -- 0x05D8
    x"FD",x"79",x"D6",x"20",x"32",x"D7",x"F3",x"3E", -- 0x05E0
    x"F1",x"C3",x"8A",x"FD",x"C5",x"D5",x"E5",x"F5", -- 0x05E8
    x"3A",x"D4",x"F3",x"C3",x"FA",x"FD",x"3A",x"D7", -- 0x05F0
    x"F3",x"3C",x"FE",x"19",x"D2",x"FF",x"FC",x"6F", -- 0x05F8
    x"CD",x"6A",x"FD",x"4F",x"3A",x"CF",x"F3",x"67", -- 0x0600
    x"3A",x"D0",x"F3",x"47",x"25",x"24",x"69",x"3A", -- 0x0608
    x"D3",x"F3",x"77",x"2C",x"C2",x"12",x"FE",x"05", -- 0x0610
    x"C2",x"0D",x"FE",x"C3",x"FF",x"FC",x"2A",x"D6", -- 0x0618
    x"F3",x"E5",x"45",x"0E",x"20",x"CD",x"37",x"FC", -- 0x0620
    x"3E",x"04",x"80",x"47",x"C2",x"25",x"FE",x"E1", -- 0x0628
    x"C3",x"FC",x"FC",x"0E",x"15",x"3A",x"E7",x"F3", -- 0x0630
    x"FB",x"3D",x"C2",x"38",x"FE",x"3A",x"E7",x"F3", -- 0x0638
    x"F3",x"3D",x"C2",x"40",x"FE",x"0D",x"C2",x"35", -- 0x0640
    x"FE",x"C9",x"C0",x"84",x"00",x"04",x"4A",x"60", -- 0x0648
    x"2A",x"1F",x"0A",x"1F",x"2A",x"11",x"0E",x"51", -- 0x0650
    x"0E",x"11",x"18",x"19",x"02",x"04",x"08",x"13", -- 0x0658
    x"03",x"04",x"2A",x"0C",x"15",x"12",x"0D",x"26", -- 0x0660
    x"02",x"04",x"40",x"02",x"04",x"48",x"04",x"02", -- 0x0668
    x"08",x"04",x"42",x"04",x"08",x"00",x"04",x"15", -- 0x0670
    x"0E",x"15",x"04",x"00",x"00",x"24",x"1F",x"24", -- 0x0678
    x"00",x"40",x"2C",x"04",x"08",x"40",x"1F",x"40", -- 0x0680
    x"80",x"2C",x"00",x"01",x"02",x"04",x"08",x"10", -- 0x0688
    x"00",x"0E",x"11",x"13",x"15",x"19",x"11",x"0E", -- 0x0690
    x"04",x"0C",x"64",x"0E",x"0E",x"11",x"01",x"06", -- 0x0698
    x"08",x"10",x"1F",x"1F",x"01",x"02",x"06",x"01", -- 0x06A0
    x"11",x"0E",x"02",x"06",x"0A",x"12",x"1F",x"22", -- 0x06A8
    x"1F",x"10",x"1E",x"21",x"11",x"0E",x"07",x"08", -- 0x06B0
    x"10",x"1E",x"31",x"0E",x"1F",x"01",x"02",x"04", -- 0x06B8
    x"48",x"0E",x"31",x"0E",x"31",x"0E",x"0E",x"31", -- 0x06C0
    x"0F",x"01",x"02",x"1C",x"00",x"2C",x"20",x"2C", -- 0x06C8
    x"2C",x"00",x"2C",x"04",x"08",x"02",x"04",x"08", -- 0x06D0
    x"10",x"08",x"04",x"02",x"20",x"1F",x"00",x"1F", -- 0x06D8
    x"20",x"08",x"04",x"02",x"01",x"02",x"04",x"08", -- 0x06E0
    x"0E",x"11",x"01",x"02",x"04",x"00",x"04",x"0E", -- 0x06E8
    x"11",x"13",x"15",x"17",x"10",x"0E",x"04",x"0A", -- 0x06F0
    x"31",x"1F",x"31",x"1E",x"31",x"1E",x"31",x"1E", -- 0x06F8
    x"0E",x"11",x"50",x"11",x"0E",x"1E",x"89",x"1E", -- 0x0700
    x"1F",x"30",x"1E",x"30",x"1F",x"1F",x"30",x"1E", -- 0x0708
    x"50",x"0E",x"11",x"30",x"13",x"11",x"0F",x"51", -- 0x0710
    x"1F",x"51",x"0E",x"84",x"0E",x"61",x"31",x"0E", -- 0x0718
    x"11",x"12",x"14",x"18",x"14",x"12",x"11",x"90", -- 0x0720
    x"11",x"1F",x"11",x"1B",x"35",x"51",x"31",x"19", -- 0x0728
    x"15",x"13",x"31",x"0E",x"91",x"0E",x"1E",x"31", -- 0x0730
    x"1E",x"50",x"0E",x"51",x"15",x"12",x"0D",x"1E", -- 0x0738
    x"31",x"1E",x"14",x"12",x"11",x"0E",x"11",x"10", -- 0x0740
    x"0E",x"01",x"11",x"0E",x"1F",x"A4",x"B1",x"0E", -- 0x0748
    x"51",x"2A",x"24",x"51",x"55",x"0A",x"31",x"0A", -- 0x0750
    x"04",x"0A",x"31",x"31",x"0A",x"64",x"1F",x"01", -- 0x0758
    x"02",x"0E",x"08",x"10",x"1F",x"0E",x"88",x"0E", -- 0x0760
    x"00",x"10",x"08",x"04",x"02",x"01",x"00",x"0E", -- 0x0768
    x"82",x"0E",x"0E",x"11",x"80",x"A0",x"1F",x"12", -- 0x0770
    x"35",x"1D",x"35",x"12",x"04",x"0A",x"31",x"1F", -- 0x0778
    x"31",x"1F",x"30",x"1E",x"31",x"1E",x"92",x"1F", -- 0x0780
    x"01",x"06",x"6A",x"1F",x"11",x"1F",x"30",x"1E", -- 0x0788
    x"30",x"1F",x"04",x"1F",x"35",x"1F",x"24",x"1F", -- 0x0790
    x"11",x"90",x"31",x"0A",x"04",x"0A",x"31",x"31", -- 0x0798
    x"13",x"15",x"19",x"31",x"15",x"11",x"13",x"15", -- 0x07A0
    x"19",x"31",x"11",x"12",x"14",x"18",x"14",x"12", -- 0x07A8
    x"11",x"07",x"89",x"19",x"11",x"1B",x"35",x"51", -- 0x07B0
    x"51",x"1F",x"51",x"0E",x"91",x"0E",x"1F",x"B1", -- 0x07B8
    x"0F",x"31",x"0F",x"05",x"09",x"11",x"1E",x"31", -- 0x07C0
    x"1E",x"50",x"0E",x"11",x"50",x"11",x"0E",x"1F", -- 0x07C8
    x"A4",x"51",x"0A",x"04",x"08",x"10",x"11",x"35", -- 0x07D0
    x"0E",x"35",x"11",x"1E",x"31",x"1E",x"31",x"1E", -- 0x07D8
    x"50",x"1E",x"31",x"1E",x"51",x"19",x"35",x"19", -- 0x07E0
    x"0E",x"11",x"01",x"06",x"01",x"11",x"0E",x"11", -- 0x07E8
    x"95",x"1F",x"0E",x"11",x"01",x"07",x"01",x"11", -- 0x07F0
    x"0E",x"95",x"1F",x"01",x"51",x"1F",x"41",x"52"  -- 0x07F8
  );

begin

  p_rom : process(clk)
  begin
    if rising_edge(clk) then
      data <= ROM(to_integer(unsigned(addr)));
    end if;
  end process;

end RTL;
