-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

entity rom_sdos is
  port (
    clk         : in    std_logic;
    addr        : in    std_logic_vector(12 downto 0);
    data        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of rom_sdos is

  type ROM_ARRAY is array(0 to 8191) of std_logic_vector(7 downto 0);
  constant ROM : ROM_ARRAY := (
    x"C3",x"30",x"B8",x"1F",x"1A",x"1A",x"20",x"28", -- 0x0000
    x"43",x"29",x"20",x"31",x"39",x"39",x"33",x"20", -- 0x0008
    x"4F",x"52",x"49",x"4F",x"4E",x"53",x"4F",x"46", -- 0x0010
    x"54",x"0D",x"0A",x"20",x"4F",x"52",x"44",x"4F", -- 0x0018
    x"53",x"20",x"56",x"34",x"2E",x"30",x"33",x"20", -- 0x0020
    x"32",x"32",x"31",x"30",x"39",x"33",x"07",x"00", -- 0x0028
    x"CD",x"12",x"F8",x"A7",x"C2",x"64",x"B8",x"CD", -- 0x0030
    x"1E",x"BB",x"32",x"60",x"B8",x"21",x"E7",x"BA", -- 0x0038
    x"3E",x"42",x"CD",x"A1",x"BE",x"CA",x"4E",x"B8", -- 0x0040
    x"21",x"4E",x"B8",x"C3",x"A8",x"BF",x"21",x"5F", -- 0x0048
    x"B8",x"22",x"46",x"B8",x"22",x"49",x"B8",x"21", -- 0x0050
    x"EB",x"BA",x"3E",x"41",x"C3",x"42",x"B8",x"3E", -- 0x0058
    x"41",x"CD",x"0B",x"BB",x"21",x"03",x"B8",x"E5", -- 0x0060
    x"CD",x"18",x"F8",x"E1",x"36",x"00",x"31",x"B9", -- 0x0068
    x"F3",x"CD",x"1A",x"BA",x"CD",x"14",x"BA",x"CD", -- 0x0070
    x"1E",x"BB",x"CD",x"16",x"BA",x"3E",x"3E",x"CD", -- 0x0078
    x"16",x"BA",x"21",x"04",x"B8",x"CD",x"57",x"BB", -- 0x0080
    x"06",x"00",x"CD",x"03",x"F8",x"FE",x"03",x"CA", -- 0x0088
    x"4E",x"BF",x"FE",x"08",x"C2",x"A9",x"B8",x"78", -- 0x0090
    x"A7",x"CA",x"8A",x"B8",x"E5",x"21",x"6B",x"B9", -- 0x0098
    x"CD",x"18",x"F8",x"E1",x"2B",x"05",x"C3",x"8A", -- 0x00A0
    x"B8",x"FE",x"0D",x"CA",x"C2",x"B8",x"FE",x"1F", -- 0x00A8
    x"DA",x"8A",x"B8",x"CD",x"16",x"BA",x"77",x"23", -- 0x00B0
    x"04",x"78",x"FE",x"1F",x"C2",x"8A",x"B8",x"C3", -- 0x00B8
    x"9C",x"B8",x"77",x"CD",x"1A",x"BA",x"21",x"04", -- 0x00C0
    x"B8",x"7E",x"47",x"23",x"FE",x"44",x"C2",x"DB", -- 0x00C8
    x"B8",x"7E",x"FE",x"3A",x"78",x"C2",x"F7",x"B8", -- 0x00D0
    x"C3",x"F0",x"B8",x"FE",x"42",x"CA",x"EA",x"B8", -- 0x00D8
    x"FE",x"43",x"CA",x"EA",x"B8",x"FE",x"41",x"C2", -- 0x00E0
    x"F7",x"B8",x"7E",x"FE",x"3A",x"C2",x"2C",x"B9", -- 0x00E8
    x"78",x"CD",x"0B",x"BB",x"23",x"7E",x"23",x"22", -- 0x00F0
    x"5B",x"BB",x"21",x"34",x"B9",x"E5",x"FE",x"44", -- 0x00F8
    x"CA",x"2C",x"BA",x"FE",x"0D",x"CA",x"2C",x"BA", -- 0x0100
    x"FE",x"52",x"CA",x"EC",x"BD",x"FE",x"53",x"CA", -- 0x0108
    x"6F",x"B9",x"FE",x"45",x"CA",x"9E",x"BA",x"FE", -- 0x0110
    x"54",x"CA",x"DB",x"B9",x"FE",x"46",x"CA",x"7B", -- 0x0118
    x"BA",x"E1",x"FE",x"4C",x"CA",x"A8",x"BF",x"FE", -- 0x0120
    x"20",x"CA",x"A8",x"BF",x"3E",x"3F",x"CD",x"16", -- 0x0128
    x"BA",x"C3",x"6E",x"B8",x"A7",x"CA",x"6E",x"B8", -- 0x0130
    x"21",x"53",x"B9",x"E5",x"21",x"AE",x"BA",x"3D", -- 0x0138
    x"C8",x"21",x"BA",x"BA",x"3D",x"C8",x"21",x"C6", -- 0x0140
    x"BA",x"3D",x"C8",x"21",x"D7",x"BA",x"3D",x"C8", -- 0x0148
    x"C3",x"2C",x"B9",x"CD",x"18",x"F8",x"2A",x"5B", -- 0x0150
    x"BB",x"7E",x"FE",x"20",x"CA",x"6E",x"B8",x"FE", -- 0x0158
    x"0D",x"CA",x"6E",x"B8",x"CD",x"16",x"BA",x"23", -- 0x0160
    x"C3",x"59",x"B9",x"08",x"20",x"08",x"00",x"2A", -- 0x0168
    x"5B",x"BB",x"7E",x"23",x"FE",x"20",x"C2",x"7C", -- 0x0170
    x"B9",x"22",x"82",x"B9",x"FE",x"0D",x"C2",x"72", -- 0x0178
    x"B9",x"21",x"00",x"00",x"EB",x"CD",x"A8",x"B9", -- 0x0180
    x"22",x"62",x"BB",x"DA",x"2C",x"B9",x"CD",x"A8", -- 0x0188
    x"B9",x"22",x"5F",x"BB",x"D2",x"2C",x"B9",x"EB", -- 0x0190
    x"2A",x"62",x"BB",x"7C",x"BA",x"DA",x"94",x"BC", -- 0x0198
    x"7D",x"BB",x"D2",x"2C",x"B9",x"C3",x"94",x"BC", -- 0x01A0
    x"21",x"00",x"00",x"45",x"4D",x"1A",x"13",x"FE", -- 0x01A8
    x"0D",x"CA",x"D9",x"B9",x"FE",x"2C",x"C8",x"D6", -- 0x01B0
    x"30",x"FA",x"2C",x"B9",x"FE",x"0A",x"FA",x"CD", -- 0x01B8
    x"B9",x"FE",x"11",x"FA",x"2C",x"B9",x"FE",x"17", -- 0x01C0
    x"F2",x"2C",x"B9",x"D6",x"07",x"4F",x"29",x"29", -- 0x01C8
    x"29",x"29",x"DA",x"2C",x"B9",x"09",x"C3",x"AD", -- 0x01D0
    x"B9",x"37",x"C9",x"CD",x"9A",x"BB",x"A7",x"3E", -- 0x01D8
    x"01",x"C8",x"CD",x"CD",x"BF",x"CD",x"21",x"BB", -- 0x01E0
    x"FE",x"0D",x"CC",x"1A",x"BA",x"E6",x"7F",x"FE", -- 0x01E8
    x"7F",x"CA",x"FF",x"B9",x"FE",x"1F",x"DA",x"FF", -- 0x01F0
    x"B9",x"CA",x"FF",x"B9",x"CD",x"16",x"BA",x"CD", -- 0x01F8
    x"1B",x"F8",x"FE",x"03",x"CA",x"28",x"BC",x"3C", -- 0x0200
    x"C2",x"FF",x"B9",x"23",x"CD",x"33",x"BD",x"C2", -- 0x0208
    x"E5",x"B9",x"AF",x"C9",x"3E",x"20",x"4F",x"C3", -- 0x0210
    x"09",x"F8",x"3E",x"0D",x"CD",x"16",x"BA",x"3E", -- 0x0218
    x"0A",x"C3",x"16",x"BA",x"7C",x"CD",x"15",x"F8", -- 0x0220
    x"7D",x"C3",x"15",x"F8",x"2A",x"9E",x"BB",x"CD", -- 0x0228
    x"14",x"BA",x"06",x"02",x"CD",x"1F",x"BC",x"A7", -- 0x0230
    x"C8",x"2A",x"03",x"BB",x"16",x"08",x"CD",x"21", -- 0x0238
    x"BB",x"CD",x"16",x"BA",x"23",x"15",x"C2",x"3E", -- 0x0240
    x"BA",x"CD",x"14",x"BA",x"CD",x"44",x"BC",x"EB", -- 0x0248
    x"CD",x"24",x"BA",x"EB",x"CD",x"14",x"BA",x"23", -- 0x0250
    x"CD",x"44",x"BC",x"EB",x"CD",x"24",x"BA",x"CD", -- 0x0258
    x"2A",x"BC",x"CD",x"12",x"F8",x"C2",x"12",x"BA", -- 0x0260
    x"16",x"04",x"CD",x"14",x"BA",x"15",x"C2",x"6A", -- 0x0268
    x"BA",x"05",x"C2",x"34",x"BA",x"CD",x"1A",x"BA", -- 0x0270
    x"C3",x"2F",x"BA",x"CD",x"90",x"BA",x"C0",x"21", -- 0x0278
    x"1F",x"BB",x"7E",x"FE",x"41",x"C2",x"8A",x"BA", -- 0x0280
    x"36",x"42",x"21",x"00",x"00",x"C3",x"5F",x"BE", -- 0x0288
    x"21",x"A5",x"BA",x"CD",x"18",x"F8",x"CD",x"03", -- 0x0290
    x"F8",x"FE",x"0D",x"3E",x"00",x"C9",x"CD",x"90", -- 0x0298
    x"BA",x"C0",x"C3",x"13",x"BE",x"20",x"64",x"61", -- 0x02A0
    x"3F",x"5B",x"77",x"6B",x"5D",x"00",x"20",x"6E", -- 0x02A8
    x"65",x"74",x"20",x"66",x"61",x"6A",x"6C",x"61", -- 0x02B0
    x"3A",x"00",x"20",x"70",x"6F",x"77",x"74",x"2E", -- 0x02B8
    x"66",x"61",x"6A",x"6C",x"3A",x"00",x"20",x"6D", -- 0x02C0
    x"61",x"6C",x"6F",x"20",x"64",x"69",x"73",x"6B", -- 0x02C8
    x"61",x"20",x"64",x"6C",x"71",x"3A",x"00",x"20", -- 0x02D0
    x"74",x"6F",x"6C",x"78",x"6B",x"6F",x"20",x"7E", -- 0x02D8
    x"74",x"65",x"6E",x"69",x"65",x"3A",x"00",x"45", -- 0x02E0
    x"58",x"54",x"20",x"56",x"43",x"20",x"20",x"53", -- 0x02E8
    x"45",x"54",x"55",x"50",x"2E",x"54",x"58",x"20", -- 0x02F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02F8
    x"C3",x"00",x"B8",x"00",x"00",x"00",x"00",x"00", -- 0x0300
    x"00",x"3E",x"41",x"E5",x"21",x"00",x"08",x"FE", -- 0x0308
    x"41",x"CA",x"17",x"BB",x"21",x"00",x"00",x"22", -- 0x0310
    x"9E",x"BB",x"E1",x"32",x"1F",x"BB",x"3E",x"41", -- 0x0318
    x"C9",x"CD",x"1E",x"BB",x"FE",x"41",x"C2",x"35", -- 0x0320
    x"BB",x"3E",x"90",x"32",x"03",x"F5",x"22",x"01", -- 0x0328
    x"F5",x"3A",x"00",x"F5",x"C9",x"E6",x"07",x"3D", -- 0x0330
    x"C5",x"CD",x"36",x"F8",x"79",x"C1",x"C9",x"7B", -- 0x0338
    x"CD",x"45",x"BB",x"23",x"7A",x"C5",x"4F",x"3A", -- 0x0340
    x"1F",x"BB",x"FE",x"41",x"CA",x"55",x"BB",x"E6", -- 0x0348
    x"07",x"3D",x"CD",x"39",x"F8",x"C1",x"C9",x"22", -- 0x0350
    x"5B",x"BB",x"21",x"00",x"00",x"C9",x"11",x"00", -- 0x0358
    x"00",x"21",x"00",x"00",x"C9",x"22",x"62",x"BB", -- 0x0360
    x"EB",x"22",x"5F",x"BB",x"C9",x"2A",x"03",x"BB", -- 0x0368
    x"44",x"4D",x"2A",x"07",x"BB",x"EB",x"2A",x"05", -- 0x0370
    x"BB",x"C9",x"2A",x"5B",x"BB",x"7E",x"FE",x"20", -- 0x0378
    x"C2",x"87",x"BB",x"23",x"C3",x"7D",x"BB",x"22", -- 0x0380
    x"5B",x"BB",x"44",x"4D",x"C9",x"22",x"91",x"BB", -- 0x0388
    x"21",x"FF",x"EF",x"C9",x"21",x"74",x"BF",x"CD", -- 0x0390
    x"57",x"BB",x"CD",x"7A",x"BB",x"21",x"00",x"08", -- 0x0398
    x"FE",x"0D",x"3E",x"00",x"C8",x"AF",x"32",x"A2", -- 0x03A0
    x"BF",x"CD",x"1F",x"BC",x"C8",x"16",x"08",x"2A", -- 0x03A8
    x"5B",x"BB",x"44",x"4D",x"2A",x"03",x"BB",x"0A", -- 0x03B0
    x"5F",x"FE",x"0D",x"CA",x"E0",x"BB",x"FE",x"20", -- 0x03B8
    x"CA",x"E0",x"BB",x"FE",x"24",x"CA",x"E0",x"BB", -- 0x03C0
    x"CD",x"21",x"BB",x"FE",x"24",x"C2",x"D3",x"BB", -- 0x03C8
    x"32",x"A2",x"BF",x"BB",x"C2",x"ED",x"BB",x"03", -- 0x03D0
    x"23",x"15",x"C2",x"B7",x"BB",x"C3",x"F6",x"BB", -- 0x03D8
    x"CD",x"21",x"BB",x"FE",x"20",x"CA",x"F6",x"BB", -- 0x03E0
    x"FE",x"24",x"CA",x"F3",x"BB",x"CD",x"2A",x"BC", -- 0x03E8
    x"C3",x"A5",x"BB",x"32",x"A2",x"BF",x"2A",x"03", -- 0x03F0
    x"BB",x"E5",x"11",x"08",x"00",x"19",x"CD",x"44", -- 0x03F8
    x"BC",x"EB",x"22",x"05",x"BB",x"EB",x"23",x"CD", -- 0x0400
    x"44",x"BC",x"23",x"23",x"23",x"23",x"23",x"22", -- 0x0408
    x"62",x"BB",x"EB",x"22",x"07",x"BB",x"19",x"22", -- 0x0410
    x"5F",x"BB",x"E1",x"3E",x"FF",x"A7",x"C9",x"22", -- 0x0418
    x"03",x"BB",x"CD",x"21",x"BB",x"FE",x"FF",x"C0", -- 0x0420
    x"AF",x"C9",x"2A",x"03",x"BB",x"E5",x"11",x"0A", -- 0x0428
    x"00",x"19",x"CD",x"44",x"BC",x"E1",x"19",x"11", -- 0x0430
    x"10",x"00",x"19",x"3E",x"00",x"17",x"A7",x"C8", -- 0x0438
    x"33",x"33",x"AF",x"C9",x"CD",x"21",x"BB",x"5F", -- 0x0440
    x"23",x"CD",x"21",x"BB",x"57",x"C9",x"C5",x"D5", -- 0x0448
    x"E5",x"CD",x"9A",x"BB",x"A7",x"C1",x"3E",x"01", -- 0x0450
    x"CA",x"74",x"BC",x"11",x"08",x"00",x"2A",x"03", -- 0x0458
    x"BB",x"19",x"CD",x"21",x"BB",x"5F",x"79",x"CD", -- 0x0460
    x"45",x"BB",x"23",x"CD",x"21",x"BB",x"57",x"78", -- 0x0468
    x"CD",x"45",x"BB",x"EB",x"D1",x"C1",x"C9",x"CD", -- 0x0470
    x"9A",x"BB",x"A7",x"3E",x"02",x"C0",x"CD",x"7A", -- 0x0478
    x"BB",x"FE",x"0D",x"CA",x"00",x"BB",x"2A",x"03", -- 0x0480
    x"BB",x"CD",x"11",x"BD",x"EB",x"2A",x"62",x"BB", -- 0x0488
    x"EB",x"C3",x"3F",x"BB",x"CD",x"77",x"BC",x"A7", -- 0x0490
    x"C0",x"23",x"E5",x"2A",x"5F",x"BB",x"EB",x"2A", -- 0x0498
    x"62",x"BB",x"7B",x"95",x"6F",x"7A",x"9C",x"67", -- 0x04A0
    x"7D",x"F6",x"0F",x"6F",x"23",x"22",x"05",x"BB", -- 0x04A8
    x"EB",x"E1",x"CD",x"3F",x"BB",x"23",x"AF",x"CD", -- 0x04B0
    x"45",x"BB",x"23",x"23",x"23",x"23",x"EB",x"21", -- 0x04B8
    x"FF",x"EF",x"3A",x"1F",x"BB",x"FE",x"42",x"C2", -- 0x04C0
    x"CD",x"BC",x"CD",x"90",x"BB",x"CD",x"33",x"BD", -- 0x04C8
    x"DA",x"07",x"BD",x"EB",x"E5",x"E5",x"2A",x"62", -- 0x04D0
    x"BB",x"4D",x"44",x"2A",x"05",x"BB",x"EB",x"E1", -- 0x04D8
    x"19",x"EB",x"E1",x"0A",x"CD",x"45",x"BB",x"23", -- 0x04E0
    x"03",x"CD",x"33",x"BD",x"CA",x"5F",x"BE",x"EB", -- 0x04E8
    x"E5",x"21",x"FF",x"EF",x"3A",x"1F",x"BB",x"FE", -- 0x04F0
    x"42",x"C2",x"FF",x"BC",x"CD",x"90",x"BB",x"CD", -- 0x04F8
    x"33",x"BD",x"E1",x"EB",x"C2",x"E3",x"BC",x"2A", -- 0x0500
    x"03",x"BB",x"CD",x"5F",x"BE",x"3E",x"03",x"A7", -- 0x0508
    x"C9",x"16",x"08",x"0A",x"FE",x"20",x"CA",x"28", -- 0x0510
    x"BD",x"FE",x"0D",x"CA",x"28",x"BD",x"CD",x"45", -- 0x0518
    x"BB",x"23",x"03",x"15",x"C2",x"13",x"BD",x"C9", -- 0x0520
    x"3E",x"20",x"CD",x"45",x"BB",x"23",x"15",x"C2", -- 0x0528
    x"28",x"BD",x"C9",x"7C",x"BA",x"C0",x"7D",x"BB", -- 0x0530
    x"C9",x"E5",x"D5",x"C5",x"C3",x"3F",x"BD",x"22", -- 0x0538
    x"62",x"BB",x"32",x"7E",x"BD",x"CD",x"77",x"BC", -- 0x0540
    x"A7",x"C2",x"C0",x"BD",x"23",x"23",x"23",x"CD", -- 0x0548
    x"45",x"BB",x"11",x"10",x"00",x"2A",x"03",x"BB", -- 0x0550
    x"19",x"22",x"AD",x"BD",x"EB",x"21",x"FF",x"EF", -- 0x0558
    x"3A",x"1F",x"BB",x"FE",x"42",x"C2",x"6B",x"BD", -- 0x0560
    x"CD",x"90",x"BB",x"CD",x"33",x"BD",x"DA",x"B7", -- 0x0568
    x"BD",x"21",x"00",x"00",x"22",x"A6",x"BD",x"21", -- 0x0570
    x"7F",x"BD",x"22",x"3D",x"BD",x"3E",x"00",x"32", -- 0x0578
    x"7E",x"BD",x"21",x"FF",x"EF",x"3A",x"1F",x"BB", -- 0x0580
    x"FE",x"42",x"C2",x"90",x"BD",x"CD",x"90",x"BB", -- 0x0588
    x"7D",x"E6",x"F0",x"6F",x"2B",x"EB",x"2A",x"AD", -- 0x0590
    x"BD",x"CD",x"33",x"BD",x"CA",x"B7",x"BD",x"3A", -- 0x0598
    x"7E",x"BD",x"CD",x"45",x"BB",x"21",x"00",x"00", -- 0x05A0
    x"23",x"22",x"A6",x"BD",x"21",x"00",x"00",x"23", -- 0x05A8
    x"22",x"AD",x"BD",x"AF",x"C3",x"C0",x"BD",x"CD", -- 0x05B0
    x"07",x"BD",x"21",x"3F",x"BD",x"22",x"3D",x"BD", -- 0x05B8
    x"C1",x"D1",x"E1",x"C9",x"21",x"3F",x"BD",x"22", -- 0x05C0
    x"3D",x"BD",x"11",x"0A",x"00",x"2A",x"03",x"BB", -- 0x05C8
    x"E5",x"19",x"EB",x"2A",x"A6",x"BD",x"2B",x"23", -- 0x05D0
    x"7D",x"E6",x"0F",x"C2",x"D7",x"BD",x"EB",x"CD", -- 0x05D8
    x"3F",x"BB",x"E1",x"19",x"11",x"10",x"00",x"19", -- 0x05E0
    x"CD",x"5F",x"BE",x"C9",x"CD",x"9A",x"BB",x"A7", -- 0x05E8
    x"3E",x"02",x"C0",x"2A",x"5B",x"BB",x"E5",x"7E", -- 0x05F0
    x"FE",x"20",x"22",x"5B",x"BB",x"23",x"C2",x"F7", -- 0x05F8
    x"BD",x"CD",x"9A",x"BB",x"A7",x"3E",x"01",x"E1", -- 0x0600
    x"C8",x"44",x"4D",x"2A",x"03",x"BB",x"CD",x"11", -- 0x0608
    x"BD",x"AF",x"C9",x"CD",x"9A",x"BB",x"3E",x"01", -- 0x0610
    x"C8",x"2A",x"03",x"BB",x"22",x"62",x"BB",x"11", -- 0x0618
    x"0C",x"00",x"19",x"CD",x"21",x"BB",x"E6",x"80", -- 0x0620
    x"3E",x"04",x"C0",x"2A",x"9E",x"BB",x"CD",x"1F", -- 0x0628
    x"BC",x"A7",x"CA",x"3B",x"BE",x"CD",x"2A",x"BC", -- 0x0630
    x"C3",x"2E",x"BE",x"2A",x"03",x"BB",x"E5",x"2A", -- 0x0638
    x"62",x"BB",x"44",x"4D",x"2A",x"5F",x"BB",x"D1", -- 0x0640
    x"CD",x"33",x"BD",x"CA",x"5D",x"BE",x"CD",x"21", -- 0x0648
    x"BB",x"E5",x"60",x"69",x"CD",x"45",x"BB",x"E1", -- 0x0650
    x"23",x"03",x"C3",x"48",x"BE",x"60",x"69",x"3E", -- 0x0658
    x"FF",x"CD",x"45",x"BB",x"C9",x"44",x"4D",x"AF", -- 0x0660
    x"32",x"93",x"BE",x"2A",x"9E",x"BB",x"CD",x"1F", -- 0x0668
    x"BC",x"A7",x"3A",x"93",x"BE",x"C8",x"2A",x"03", -- 0x0670
    x"BB",x"E5",x"11",x"0C",x"00",x"19",x"CD",x"21", -- 0x0678
    x"BB",x"E1",x"0F",x"DA",x"98",x"BE",x"16",x"10", -- 0x0680
    x"CD",x"21",x"BB",x"02",x"23",x"03",x"15",x"C2", -- 0x0688
    x"88",x"BE",x"3E",x"00",x"3C",x"32",x"93",x"BE", -- 0x0690
    x"CD",x"2A",x"BC",x"C3",x"6E",x"BE",x"21",x"EF", -- 0x0698
    x"BA",x"CD",x"0B",x"BB",x"CD",x"57",x"BB",x"C3", -- 0x06A0
    x"9A",x"BB",x"31",x"B9",x"F3",x"CD",x"12",x"F8", -- 0x06A8
    x"A7",x"C2",x"00",x"BB",x"21",x"00",x"00",x"06", -- 0x06B0
    x"03",x"3E",x"01",x"CD",x"36",x"F8",x"79",x"FE", -- 0x06B8
    x"20",x"DA",x"D1",x"BE",x"FE",x"7F",x"D2",x"D1", -- 0x06C0
    x"BE",x"23",x"05",x"C2",x"B9",x"BE",x"C3",x"DC", -- 0x06C8
    x"BE",x"21",x"00",x"00",x"3A",x"BA",x"BE",x"0E", -- 0x06D0
    x"FF",x"CD",x"39",x"F8",x"3A",x"BA",x"BE",x"3C", -- 0x06D8
    x"FE",x"04",x"32",x"BA",x"BE",x"C2",x"B4",x"BE", -- 0x06E0
    x"3E",x"42",x"CD",x"9E",x"BE",x"C2",x"F8",x"BE", -- 0x06E8
    x"3E",x"41",x"CD",x"9E",x"BE",x"CA",x"3F",x"BF", -- 0x06F0
    x"21",x"4E",x"BF",x"22",x"FE",x"BF",x"21",x"04", -- 0x06F8
    x"BF",x"C3",x"A8",x"BF",x"EB",x"22",x"0C",x"BF", -- 0x0700
    x"31",x"B9",x"F3",x"21",x"00",x"00",x"7E",x"FE", -- 0x0708
    x"2E",x"CA",x"3F",x"BF",x"4F",x"CD",x"57",x"BB", -- 0x0710
    x"23",x"7E",x"FE",x"3A",x"C2",x"27",x"BF",x"23", -- 0x0718
    x"CD",x"57",x"BB",x"79",x"CD",x"0B",x"BB",x"7E", -- 0x0720
    x"FE",x"2E",x"CA",x"33",x"BF",x"23",x"FE",x"0D", -- 0x0728
    x"C2",x"27",x"BF",x"22",x"0C",x"BF",x"21",x"08", -- 0x0730
    x"BF",x"22",x"FE",x"BF",x"C3",x"A8",x"BF",x"21", -- 0x0738
    x"FF",x"BA",x"CD",x"33",x"F8",x"21",x"4E",x"BF", -- 0x0740
    x"22",x"FE",x"BF",x"CD",x"09",x"BB",x"31",x"B9", -- 0x0748
    x"F3",x"3A",x"1F",x"BB",x"F5",x"CD",x"09",x"BB", -- 0x0750
    x"01",x"00",x"B8",x"21",x"00",x"00",x"11",x"03", -- 0x0758
    x"03",x"CD",x"21",x"BB",x"02",x"03",x"23",x"1B", -- 0x0760
    x"7B",x"B2",x"C2",x"61",x"BF",x"F1",x"CD",x"0B", -- 0x0768
    x"BB",x"C3",x"00",x"BB",x"3F",x"26",x"20",x"00", -- 0x0770
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0778
    x"CD",x"9A",x"BB",x"A7",x"3E",x"01",x"C8",x"2A", -- 0x0780
    x"05",x"BB",x"22",x"9F",x"BF",x"44",x"4D",x"CD", -- 0x0788
    x"5E",x"BB",x"CD",x"21",x"BB",x"02",x"23",x"03", -- 0x0790
    x"CD",x"33",x"BD",x"C2",x"92",x"BF",x"21",x"00", -- 0x0798
    x"00",x"3E",x"00",x"A7",x"C8",x"3E",x"80",x"C9", -- 0x07A0
    x"22",x"B0",x"BF",x"CD",x"80",x"BF",x"EB",x"21", -- 0x07A8
    x"FD",x"BF",x"E5",x"FE",x"80",x"C0",x"EB",x"E9", -- 0x07B0
    x"C3",x"94",x"BB",x"3E",x"40",x"C9",x"C3",x"4E", -- 0x07B8
    x"BC",x"C3",x"90",x"BB",x"C3",x"8D",x"BB",x"C3", -- 0x07C0
    x"6D",x"BB",x"C3",x"65",x"BB",x"C3",x"5E",x"BB", -- 0x07C8
    x"C3",x"57",x"BB",x"C3",x"5A",x"BB",x"C3",x"0B", -- 0x07D0
    x"BB",x"C3",x"1E",x"BB",x"C3",x"21",x"BB",x"C3", -- 0x07D8
    x"45",x"BB",x"C3",x"5F",x"BE",x"C3",x"9A",x"BB", -- 0x07E0
    x"C3",x"65",x"BE",x"C3",x"EC",x"BD",x"C3",x"13", -- 0x07E8
    x"BE",x"C3",x"39",x"BD",x"C3",x"C4",x"BD",x"C3", -- 0x07F0
    x"94",x"BC",x"C3",x"80",x"BF",x"C3",x"AA",x"BE", -- 0x07F8
    x"56",x"43",x"24",x"20",x"20",x"20",x"20",x"20", -- 0x0800
    x"00",x"AD",x"00",x"0E",x"00",x"FF",x"FF",x"FF", -- 0x0808
    x"C3",x"1D",x"AD",x"C3",x"93",x"AD",x"00",x"00", -- 0x0810
    x"00",x"41",x"42",x"43",x"44",x"00",x"00",x"00", -- 0x0818
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0820
    x"00",x"00",x"00",x"00",x"FF",x"31",x"C0",x"F3", -- 0x0828
    x"CD",x"62",x"AF",x"3A",x"87",x"F3",x"E6",x"C0", -- 0x0830
    x"CA",x"37",x"AD",x"31",x"C0",x"F3",x"21",x"72", -- 0x0838
    x"F3",x"11",x"06",x"AD",x"CD",x"6D",x"B7",x"21", -- 0x0840
    x"00",x"AD",x"22",x"01",x"BB",x"CD",x"EB",x"B3", -- 0x0848
    x"21",x"00",x"F3",x"11",x"0C",x"B8",x"CD",x"6D", -- 0x0850
    x"B7",x"2B",x"11",x"02",x"B8",x"CD",x"6D",x"B7", -- 0x0858
    x"CD",x"61",x"B6",x"CD",x"03",x"F3",x"CD",x"53", -- 0x0860
    x"B3",x"CD",x"4C",x"B3",x"11",x"FF",x"FF",x"1C", -- 0x0868
    x"CD",x"3E",x"AE",x"CA",x"5F",x"AD",x"14",x"CD", -- 0x0870
    x"19",x"B0",x"CD",x"FC",x"AD",x"CA",x"66",x"AD", -- 0x0878
    x"7A",x"93",x"5F",x"1C",x"1D",x"CA",x"7E",x"AD", -- 0x0880
    x"CD",x"3E",x"AE",x"C3",x"74",x"AD",x"CD",x"C2", -- 0x0888
    x"B4",x"C3",x"93",x"AD",x"CD",x"EB",x"B3",x"CD", -- 0x0890
    x"61",x"B6",x"CD",x"C2",x"B4",x"31",x"C0",x"F3", -- 0x0898
    x"CD",x"E7",x"AF",x"21",x"93",x"AD",x"E5",x"CD", -- 0x08A0
    x"5C",x"AF",x"CD",x"71",x"B0",x"FE",x"40",x"DA", -- 0x08A8
    x"A4",x"AD",x"E6",x"5F",x"F5",x"CD",x"EC",x"AD", -- 0x08B0
    x"F1",x"FE",x"4D",x"CA",x"96",x"AE",x"FE",x"58", -- 0x08B8
    x"CA",x"93",x"AE",x"FE",x"0D",x"C2",x"C3",x"AD", -- 0x08C0
    x"3A",x"7D",x"F3",x"47",x"B7",x"CA",x"84",x"AE", -- 0x08C8
    x"C3",x"F2",x"B7",x"FE",x"53",x"CA",x"BA",x"B9", -- 0x08D0
    x"4F",x"AF",x"B0",x"C8",x"79",x"FE",x"45",x"CA", -- 0x08D8
    x"4B",x"B8",x"FE",x"43",x"CA",x"CC",x"B8",x"FE", -- 0x08E0
    x"52",x"CA",x"5F",x"B5",x"FE",x"4C",x"CA",x"DE", -- 0x08E8
    x"B7",x"FE",x"54",x"CA",x"B8",x"BA",x"FE",x"41", -- 0x08F0
    x"CA",x"FF",x"AE",x"C9",x"FE",x"03",x"CA",x"00", -- 0x08F8
    x"AD",x"FE",x"18",x"CA",x"FC",x"AD",x"FE",x"08", -- 0x0900
    x"CA",x"3E",x"AE",x"C9",x"CD",x"81",x"AF",x"CA", -- 0x0908
    x"14",x"AE",x"E6",x"04",x"79",x"C0",x"E6",x"01", -- 0x0910
    x"79",x"CA",x"0D",x"AE",x"C9",x"3C",x"32",x"87", -- 0x0918
    x"F3",x"C3",x"2D",x"AE",x"E6",x"10",x"79",x"C2", -- 0x0920
    x"27",x"AE",x"E6",x"01",x"79",x"CA",x"0D",x"AE", -- 0x0928
    x"E6",x"FC",x"F6",x"02",x"C3",x"0E",x"AE",x"CD", -- 0x0930
    x"20",x"AE",x"C3",x"2D",x"AE",x"E5",x"21",x"72", -- 0x0938
    x"F3",x"0E",x"12",x"23",x"7E",x"2B",x"77",x"23", -- 0x0940
    x"0D",x"C2",x"33",x"AE",x"E1",x"C9",x"CD",x"81", -- 0x0948
    x"AF",x"CA",x"63",x"AE",x"E6",x"04",x"79",x"C2", -- 0x0950
    x"50",x"AE",x"E6",x"01",x"79",x"C2",x"6F",x"AE", -- 0x0958
    x"E6",x"FC",x"4F",x"E6",x"10",x"79",x"CA",x"5F", -- 0x0960
    x"AE",x"CD",x"70",x"AE",x"C3",x"73",x"AE",x"3C", -- 0x0968
    x"C3",x"70",x"AE",x"E6",x"10",x"79",x"C0",x"E6", -- 0x0970
    x"01",x"79",x"C2",x"6F",x"AE",x"3C",x"C9",x"3D", -- 0x0978
    x"32",x"87",x"F3",x"E5",x"21",x"84",x"F3",x"0E", -- 0x0980
    x"12",x"2B",x"7E",x"23",x"77",x"2B",x"0D",x"C2", -- 0x0988
    x"79",x"AE",x"E1",x"C9",x"21",x"8D",x"AD",x"E5", -- 0x0990
    x"21",x"75",x"F3",x"34",x"7E",x"FE",x"45",x"C0", -- 0x0998
    x"36",x"41",x"C9",x"CD",x"9A",x"AE",x"21",x"8D", -- 0x09A0
    x"AD",x"E5",x"CD",x"81",x"AF",x"11",x"30",x"10", -- 0x09A8
    x"21",x"85",x"F3",x"CA",x"AA",x"AE",x"11",x"0C", -- 0x09B0
    x"04",x"23",x"A3",x"C2",x"C2",x"AE",x"79",x"E6", -- 0x09B8
    x"01",x"CA",x"BA",x"AE",x"CD",x"3E",x"AE",x"CD", -- 0x09C0
    x"DE",x"AE",x"3A",x"87",x"F3",x"82",x"32",x"87", -- 0x09C8
    x"F3",x"C9",x"82",x"A3",x"CA",x"C8",x"AE",x"82", -- 0x09D0
    x"F5",x"F5",x"7B",x"2F",x"A1",x"4F",x"F1",x"B1", -- 0x09D8
    x"32",x"87",x"F3",x"F1",x"C0",x"7E",x"3C",x"C0", -- 0x09E0
    x"CD",x"DE",x"AE",x"C3",x"FC",x"AD",x"E5",x"D5", -- 0x09E8
    x"7E",x"2F",x"77",x"21",x"75",x"F3",x"06",x"04", -- 0x09F0
    x"23",x"5E",x"2B",x"7E",x"73",x"23",x"77",x"23", -- 0x09F8
    x"23",x"23",x"05",x"C2",x"E8",x"AE",x"D1",x"E1", -- 0x0A00
    x"C9",x"CD",x"55",x"BA",x"C3",x"17",x"AF",x"CD", -- 0x0A08
    x"70",x"AF",x"FE",x"01",x"CA",x"17",x"AF",x"C9", -- 0x0A10
    x"F5",x"CD",x"9A",x"AE",x"F1",x"B7",x"C4",x"9A", -- 0x0A18
    x"AE",x"CD",x"E7",x"AF",x"CD",x"E5",x"B1",x"2A", -- 0x0A20
    x"4C",x"F3",x"7D",x"C6",x"0A",x"6F",x"CD",x"3C", -- 0x0A28
    x"F8",x"21",x"53",x"AF",x"CD",x"18",x"F8",x"0E", -- 0x0A30
    x"05",x"CD",x"16",x"B6",x"36",x"0D",x"11",x"5A", -- 0x0A38
    x"F3",x"CD",x"70",x"BA",x"C2",x"F9",x"AE",x"D2", -- 0x0A40
    x"F9",x"AE",x"EB",x"D5",x"2A",x"4A",x"F3",x"E5", -- 0x0A48
    x"CD",x"D0",x"BF",x"EB",x"CD",x"BE",x"BF",x"E1", -- 0x0A50
    x"3E",x"08",x"85",x"6F",x"D1",x"73",x"23",x"72", -- 0x0A58
    x"C3",x"3D",x"B7",x"20",x"20",x"20",x"20",x"08", -- 0x0A60
    x"08",x"08",x"08",x"00",x"CD",x"62",x"AF",x"C3", -- 0x0A68
    x"D6",x"BF",x"3A",x"75",x"F3",x"FE",x"41",x"DA", -- 0x0A70
    x"2B",x"AD",x"FE",x"45",x"D2",x"2B",x"AD",x"C9", -- 0x0A78
    x"C5",x"CD",x"81",x"AF",x"C2",x"79",x"AF",x"0F", -- 0x0A80
    x"0F",x"E6",x"0C",x"0F",x"0F",x"FE",x"03",x"C1", -- 0x0A88
    x"C9",x"3A",x"87",x"F3",x"4F",x"E6",x"02",x"79", -- 0x0A90
    x"C9",x"CD",x"62",x"AF",x"CD",x"E4",x"B6",x"78", -- 0x0A98
    x"3C",x"32",x"81",x"F3",x"C5",x"3A",x"79",x"F3", -- 0x0AA0
    x"B8",x"DA",x"A0",x"AF",x"AF",x"32",x"79",x"F3", -- 0x0AA8
    x"F5",x"22",x"3B",x"B2",x"CD",x"24",x"B3",x"7C", -- 0x0AB0
    x"32",x"97",x"B2",x"32",x"E6",x"B2",x"78",x"32", -- 0x0AB8
    x"92",x"B2",x"32",x"E1",x"B2",x"3E",x"0A",x"32", -- 0x0AC0
    x"99",x"B2",x"CD",x"70",x"AF",x"3E",x"13",x"32", -- 0x0AC8
    x"A3",x"B2",x"C2",x"C6",x"AF",x"87",x"32",x"8F", -- 0x0AD0
    x"B1",x"32",x"04",x"B2",x"32",x"56",x"B0",x"47", -- 0x0AD8
    x"F1",x"80",x"4F",x"3A",x"7D",x"F3",x"B9",x"DA", -- 0x0AE0
    x"E0",x"AF",x"3A",x"79",x"F3",x"32",x"7D",x"F3", -- 0x0AE8
    x"C1",x"B8",x"D8",x"78",x"C3",x"1D",x"B1",x"CD", -- 0x0AF0
    x"81",x"AF",x"21",x"4C",x"B3",x"06",x"0C",x"C2", -- 0x0AF8
    x"F7",x"AF",x"21",x"53",x"B3",x"06",x"30",x"C5", -- 0x0B00
    x"F5",x"11",x"FE",x"AF",x"D5",x"E9",x"F1",x"C1", -- 0x0B08
    x"A0",x"79",x"C2",x"19",x"B0",x"E6",x"01",x"CA", -- 0x0B10
    x"13",x"B0",x"CD",x"16",x"B0",x"CD",x"FC",x"AD", -- 0x0B18
    x"C3",x"19",x"B0",x"CD",x"0D",x"B0",x"CD",x"3E", -- 0x0B20
    x"AE",x"D5",x"F5",x"CD",x"C8",x"B1",x"2C",x"2C", -- 0x0B28
    x"26",x"00",x"CD",x"3C",x"F8",x"CD",x"61",x"B2", -- 0x0B30
    x"CD",x"62",x"AF",x"CD",x"0F",x"F8",x"3E",x"3A", -- 0x0B38
    x"CD",x"0F",x"F8",x"2D",x"2D",x"CD",x"72",x"B6", -- 0x0B40
    x"3A",x"7D",x"F3",x"F5",x"3A",x"79",x"F3",x"4F", -- 0x0B48
    x"CD",x"70",x"AF",x"79",x"C2",x"55",x"B0",x"E6", -- 0x0B50
    x"01",x"79",x"CA",x"55",x"B0",x"3D",x"32",x"79", -- 0x0B58
    x"F3",x"21",x"7D",x"F3",x"35",x"06",x"00",x"CD", -- 0x0B60
    x"E2",x"B1",x"05",x"CA",x"6A",x"B0",x"3A",x"81", -- 0x0B68
    x"F3",x"4F",x"3A",x"7D",x"F3",x"3C",x"B9",x"DA", -- 0x0B70
    x"57",x"B0",x"F1",x"32",x"7D",x"F3",x"F1",x"D1", -- 0x0B78
    x"C9",x"CD",x"89",x"AF",x"CD",x"7F",x"B2",x"11", -- 0x0B80
    x"74",x"B0",x"D5",x"CD",x"0A",x"B7",x"F5",x"CD", -- 0x0B88
    x"E5",x"B1",x"F1",x"FE",x"00",x"CA",x"E3",x"B0", -- 0x0B90
    x"FE",x"02",x"CA",x"A8",x"B0",x"FE",x"1A",x"CA", -- 0x0B98
    x"70",x"B1",x"FE",x"19",x"CA",x"05",x"B1",x"FE", -- 0x0BA0
    x"08",x"CA",x"AB",x"B1",x"FE",x"18",x"CA",x"97", -- 0x0BA8
    x"B1",x"FE",x"0C",x"CA",x"BF",x"B1",x"E1",x"C9", -- 0x0BB0
    x"3A",x"79",x"F3",x"4F",x"3A",x"7D",x"F3",x"91", -- 0x0BB8
    x"47",x"CD",x"70",x"AF",x"79",x"C2",x"BA",x"B0", -- 0x0BC0
    x"C6",x"12",x"C6",x"12",x"4F",x"3A",x"81",x"F3", -- 0x0BC8
    x"3D",x"B9",x"D8",x"79",x"32",x"7D",x"F3",x"0E", -- 0x0BD0
    x"0A",x"C5",x"CD",x"70",x"B1",x"CD",x"E5",x"B1", -- 0x0BD8
    x"C1",x"0D",x"C2",x"C9",x"B0",x"3A",x"81",x"F3", -- 0x0BE0
    x"4F",x"3A",x"79",x"F3",x"80",x"91",x"D0",x"81", -- 0x0BE8
    x"C3",x"1D",x"B1",x"3A",x"79",x"F3",x"4F",x"3A", -- 0x0BF0
    x"7D",x"F3",x"91",x"47",x"79",x"32",x"7D",x"F3", -- 0x0BF8
    x"0E",x"0A",x"C5",x"CD",x"05",x"B1",x"CD",x"E5", -- 0x0C00
    x"B1",x"C1",x"0D",x"C2",x"F2",x"B0",x"3A",x"79", -- 0x0C08
    x"F3",x"80",x"C3",x"1D",x"B1",x"CD",x"70",x"AF", -- 0x0C10
    x"3E",x"01",x"C2",x"0E",x"B1",x"3C",x"47",x"3A", -- 0x0C18
    x"79",x"F3",x"4F",x"3A",x"7D",x"F3",x"90",x"D8", -- 0x0C20
    x"91",x"DA",x"21",x"B1",x"81",x"32",x"7D",x"F3", -- 0x0C28
    x"C9",x"81",x"F5",x"CD",x"70",x"AF",x"3E",x"01", -- 0x0C30
    x"C2",x"2C",x"B1",x"3C",x"4F",x"3A",x"79",x"F3", -- 0x0C38
    x"91",x"32",x"79",x"F3",x"CD",x"D9",x"B2",x"F1", -- 0x0C40
    x"4F",x"CD",x"70",x"AF",x"79",x"C2",x"1D",x"B1", -- 0x0C48
    x"E6",x"01",x"CA",x"4D",x"B1",x"0D",x"CD",x"E1", -- 0x0C50
    x"B1",x"0C",x"C3",x"52",x"B1",x"0C",x"CD",x"E1", -- 0x0C58
    x"B1",x"0D",x"79",x"C3",x"1D",x"B1",x"81",x"F5", -- 0x0C60
    x"CD",x"70",x"AF",x"3E",x"01",x"C2",x"61",x"B1", -- 0x0C68
    x"3C",x"4F",x"3A",x"79",x"F3",x"81",x"32",x"79", -- 0x0C70
    x"F3",x"CD",x"8A",x"B2",x"F1",x"C3",x"38",x"B1", -- 0x0C78
    x"CD",x"70",x"AF",x"3E",x"01",x"C2",x"79",x"B1", -- 0x0C80
    x"3C",x"47",x"3A",x"7D",x"F3",x"80",x"4F",x"3A", -- 0x0C88
    x"81",x"F3",x"3D",x"B9",x"D8",x"3A",x"79",x"F3", -- 0x0C90
    x"4F",x"3A",x"7D",x"F3",x"91",x"80",x"FE",x"00", -- 0x0C98
    x"D2",x"56",x"B1",x"81",x"C3",x"1D",x"B1",x"CD", -- 0x0CA0
    x"70",x"AF",x"06",x"01",x"C2",x"A7",x"B1",x"3A", -- 0x0CA8
    x"7D",x"F3",x"E6",x"01",x"CA",x"7A",x"B1",x"E1", -- 0x0CB0
    x"3E",x"18",x"C9",x"CD",x"70",x"AF",x"06",x"01", -- 0x0CB8
    x"C2",x"BB",x"B1",x"3A",x"7D",x"F3",x"E6",x"01", -- 0x0CC0
    x"C2",x"0F",x"B1",x"E1",x"3E",x"08",x"C9",x"3A", -- 0x0CC8
    x"79",x"F3",x"32",x"7D",x"F3",x"C3",x"1D",x"B1", -- 0x0CD0
    x"3A",x"87",x"F3",x"E6",x"03",x"4F",x"CD",x"70", -- 0x0CD8
    x"AF",x"E6",x"01",x"79",x"CA",x"D9",x"B1",x"E6", -- 0x0CE0
    x"02",x"07",x"07",x"07",x"07",x"C6",x"02",x"6F", -- 0x0CE8
    x"C9",x"79",x"32",x"7D",x"F3",x"C5",x"CD",x"EB", -- 0x0CF0
    x"B1",x"C1",x"C9",x"CD",x"C8",x"B1",x"26",x"02", -- 0x0CF8
    x"3A",x"81",x"F3",x"4F",x"3A",x"7D",x"F3",x"B9", -- 0x0D00
    x"D0",x"3A",x"79",x"F3",x"4F",x"3A",x"7D",x"F3", -- 0x0D08
    x"91",x"D8",x"E5",x"FE",x"00",x"E1",x"D0",x"F5", -- 0x0D10
    x"CD",x"70",x"AF",x"CA",x"13",x"B2",x"F1",x"4F", -- 0x0D18
    x"C3",x"1D",x"B2",x"F1",x"0F",x"4F",x"D2",x"1D", -- 0x0D20
    x"B2",x"7D",x"C6",x"0E",x"6F",x"79",x"E6",x"7F", -- 0x0D28
    x"84",x"67",x"22",x"4C",x"F3",x"CD",x"3C",x"F8", -- 0x0D30
    x"CD",x"61",x"B2",x"3A",x"7D",x"F3",x"B7",x"CA", -- 0x0D38
    x"66",x"B2",x"3D",x"6F",x"26",x"00",x"29",x"29", -- 0x0D40
    x"29",x"29",x"01",x"00",x"A0",x"09",x"06",x"00", -- 0x0D48
    x"22",x"4A",x"F3",x"7E",x"CD",x"0F",x"F8",x"23", -- 0x0D50
    x"04",x"78",x"FE",x"08",x"C2",x"43",x"B2",x"CD", -- 0x0D58
    x"61",x"B2",x"CD",x"70",x"AF",x"FE",x"01",x"C0", -- 0x0D60
    x"CD",x"93",x"B6",x"CD",x"61",x"B2",x"CD",x"7D", -- 0x0D68
    x"B6",x"3E",x"20",x"C3",x"0F",x"F8",x"3E",x"2E", -- 0x0D70
    x"CD",x"0F",x"F8",x"CD",x"0F",x"F8",x"CD",x"70", -- 0x0D78
    x"AF",x"0E",x"07",x"FE",x"01",x"3E",x"20",x"C2", -- 0x0D80
    x"FB",x"B5",x"0E",x"18",x"C3",x"FB",x"B5",x"CD", -- 0x0D88
    x"85",x"B2",x"CD",x"E5",x"B1",x"3E",x"7F",x"C3", -- 0x0D90
    x"0F",x"F8",x"21",x"00",x"00",x"39",x"22",x"D6", -- 0x0D98
    x"B2",x"3E",x"00",x"32",x"CD",x"B2",x"26",x"00", -- 0x0DA0
    x"3E",x"0A",x"C6",x"14",x"6F",x"F9",x"7D",x"D6", -- 0x0DA8
    x"0A",x"6F",x"3E",x"13",x"3D",x"D1",x"C1",x"73", -- 0x0DB0
    x"2C",x"72",x"2C",x"71",x"2C",x"70",x"2C",x"D1", -- 0x0DB8
    x"C1",x"73",x"2C",x"72",x"2C",x"71",x"2C",x"70", -- 0x0DC0
    x"2C",x"D1",x"73",x"2C",x"72",x"2C",x"3D",x"C2", -- 0x0DC8
    x"A5",x"B2",x"3E",x"0A",x"36",x"00",x"2C",x"3D", -- 0x0DD0
    x"C2",x"C4",x"B2",x"24",x"3E",x"00",x"3D",x"32", -- 0x0DD8
    x"CD",x"B2",x"C2",x"98",x"B2",x"31",x"00",x"00", -- 0x0DE0
    x"C9",x"21",x"00",x"00",x"39",x"22",x"D6",x"B2", -- 0x0DE8
    x"3E",x"00",x"32",x"19",x"B3",x"26",x"00",x"2E", -- 0x0DF0
    x"D2",x"F9",x"7D",x"D6",x"0A",x"6F",x"3E",x"13", -- 0x0DF8
    x"3D",x"2D",x"56",x"2D",x"5E",x"2D",x"46",x"2D", -- 0x0E00
    x"4E",x"D5",x"C5",x"2D",x"56",x"2D",x"5E",x"2D", -- 0x0E08
    x"46",x"2D",x"4E",x"D5",x"C5",x"2D",x"56",x"2D", -- 0x0E10
    x"5E",x"D5",x"3D",x"C2",x"F1",x"B2",x"3E",x"0A", -- 0x0E18
    x"36",x"00",x"2C",x"3D",x"C2",x"10",x"B3",x"24", -- 0x0E20
    x"3E",x"00",x"3D",x"32",x"19",x"B3",x"C2",x"E7", -- 0x0E28
    x"B2",x"C3",x"D5",x"B2",x"CD",x"70",x"AF",x"E6", -- 0x0E30
    x"01",x"3A",x"87",x"F3",x"26",x"C1",x"C2",x"42", -- 0x0E38
    x"B3",x"E6",x"03",x"06",x"0A",x"B7",x"C8",x"26", -- 0x0E40
    x"CC",x"3D",x"C8",x"26",x"D9",x"3D",x"C8",x"26", -- 0x0E48
    x"E4",x"C9",x"E6",x"02",x"CA",x"49",x"B3",x"26", -- 0x0E50
    x"D9",x"06",x"16",x"C9",x"26",x"D8",x"0E",x"0C", -- 0x0E58
    x"C3",x"57",x"B3",x"26",x"C0",x"0E",x"30",x"3A", -- 0x0E60
    x"87",x"F3",x"A1",x"F5",x"01",x"E6",x"17",x"2E", -- 0x0E68
    x"00",x"CD",x"6C",x"B4",x"2E",x"04",x"0E",x"E0", -- 0x0E70
    x"CD",x"8A",x"B3",x"2E",x"D8",x"06",x"16",x"36", -- 0x0E78
    x"FF",x"24",x"05",x"C2",x"6F",x"B3",x"F1",x"C0", -- 0x0E80
    x"3E",x"F4",x"84",x"67",x"0E",x"DF",x"2E",x"07", -- 0x0E88
    x"2C",x"3E",x"01",x"B6",x"77",x"0D",x"C2",x"80", -- 0x0E90
    x"B3",x"C9",x"D5",x"E5",x"C5",x"78",x"06",x"0F", -- 0x0E98
    x"E5",x"C5",x"F5",x"11",x"09",x"08",x"CD",x"B4", -- 0x0EA0
    x"B3",x"F1",x"C1",x"E1",x"84",x"67",x"11",x"90", -- 0x0EA8
    x"10",x"3E",x"01",x"06",x"F0",x"CD",x"B4",x"B3", -- 0x0EB0
    x"C1",x"E1",x"05",x"24",x"7D",x"C6",x"04",x"6F", -- 0x0EB8
    x"0D",x"0D",x"D1",x"C9",x"32",x"E0",x"B3",x"70", -- 0x0EC0
    x"CD",x"C7",x"B3",x"73",x"2C",x"0D",x"C2",x"BB", -- 0x0EC8
    x"B3",x"2D",x"CD",x"C7",x"B3",x"70",x"C9",x"C5", -- 0x0ED0
    x"CD",x"DA",x"B3",x"CD",x"D7",x"B3",x"CD",x"D7", -- 0x0ED8
    x"B3",x"2C",x"CD",x"DA",x"B3",x"C1",x"C9",x"2C", -- 0x0EE0
    x"72",x"01",x"01",x"00",x"00",x"0D",x"E5",x"3E", -- 0x0EE8
    x"00",x"46",x"70",x"41",x"24",x"3D",x"C2",x"E2", -- 0x0EF0
    x"B3",x"E1",x"C9",x"01",x"41",x"04",x"11",x"4E", -- 0x0EF8
    x"F3",x"AF",x"21",x"00",x"A0",x"E5",x"E1",x"3C", -- 0x0F00
    x"CD",x"FE",x"B6",x"E5",x"D5",x"C5",x"79",x"CD", -- 0x0F08
    x"D6",x"BF",x"CD",x"E8",x"BF",x"C1",x"D1",x"EB", -- 0x0F10
    x"77",x"23",x"73",x"23",x"72",x"23",x"0C",x"EB", -- 0x0F18
    x"05",x"C2",x"F6",x"B3",x"E1",x"C9",x"16",x"1F", -- 0x0F20
    x"01",x"16",x"9F",x"C3",x"26",x"B4",x"CD",x"3D", -- 0x0F28
    x"B7",x"16",x"1F",x"2A",x"4C",x"F3",x"CD",x"3C", -- 0x0F30
    x"F8",x"01",x"0A",x"16",x"CD",x"70",x"AF",x"FE", -- 0x0F38
    x"01",x"CA",x"36",x"B4",x"06",x"08",x"C3",x"3B", -- 0x0F40
    x"B4",x"16",x"4E",x"CD",x"1E",x"F8",x"7D",x"85", -- 0x0F48
    x"85",x"6C",x"0F",x"0F",x"E6",x"3F",x"C6",x"C0", -- 0x0F50
    x"67",x"7D",x"85",x"07",x"85",x"07",x"6F",x"C3", -- 0x0F58
    x"5F",x"B4",x"3E",x"F0",x"32",x"E9",x"D7",x"21", -- 0x0F60
    x"EA",x"C0",x"01",x"16",x"30",x"16",x"1F",x"E5", -- 0x0F68
    x"CD",x"8F",x"B4",x"E1",x"F5",x"CD",x"6E",x"B4", -- 0x0F70
    x"F1",x"CD",x"AB",x"B4",x"37",x"3F",x"E5",x"C5", -- 0x0F78
    x"E5",x"C5",x"36",x"00",x"DC",x"06",x"F3",x"2C", -- 0x0F80
    x"0D",x"C2",x"72",x"B4",x"C1",x"E1",x"24",x"05", -- 0x0F88
    x"C2",x"70",x"B4",x"C1",x"E1",x"C9",x"CD",x"5C", -- 0x0F90
    x"AF",x"21",x"8F",x"B4",x"C3",x"B8",x"B4",x"D5", -- 0x0F98
    x"C5",x"3E",x"42",x"CD",x"D6",x"BF",x"CD",x"89", -- 0x0FA0
    x"B4",x"CD",x"5C",x"AF",x"7C",x"FE",x"C0",x"C1", -- 0x0FA8
    x"D1",x"C9",x"CD",x"62",x"AF",x"FE",x"42",x"C0", -- 0x0FB0
    x"7C",x"FE",x"C0",x"3E",x"07",x"DA",x"B1",x"B4", -- 0x0FB8
    x"AF",x"32",x"00",x"F8",x"C9",x"2A",x"4A",x"F3", -- 0x0FC0
    x"CD",x"D0",x"BF",x"C3",x"E5",x"BF",x"18",x"20", -- 0x0FC8
    x"20",x"00",x"CD",x"52",x"B4",x"21",x"36",x"B5", -- 0x0FD0
    x"E5",x"21",x"02",x"18",x"CD",x"3C",x"F8",x"01", -- 0x0FD8
    x"0C",x"02",x"16",x"0E",x"CD",x"3B",x"B4",x"E1", -- 0x0FE0
    x"7E",x"23",x"E5",x"21",x"BF",x"B4",x"77",x"2B", -- 0x0FE8
    x"CD",x"18",x"F8",x"CD",x"1E",x"F8",x"7D",x"C6", -- 0x0FF0
    x"05",x"FE",x"3F",x"6F",x"DA",x"CC",x"B4",x"CD", -- 0x0FF8
    x"1F",x"B5",x"AF",x"32",x"29",x"B5",x"CD",x"1F", -- 0x1000
    x"B5",x"CD",x"1F",x"B5",x"3E",x"B6",x"32",x"29", -- 0x1008
    x"B5",x"21",x"04",x"18",x"D1",x"06",x"03",x"E5", -- 0x1010
    x"CD",x"3C",x"F8",x"1A",x"CD",x"0F",x"F8",x"13", -- 0x1018
    x"05",x"C2",x"0B",x"B5",x"E1",x"7D",x"C6",x"08", -- 0x1020
    x"6F",x"FE",x"3F",x"DA",x"05",x"B5",x"C9",x"2E", -- 0x1028
    x"F0",x"26",x"EF",x"06",x"30",x"AF",x"7E",x"17", -- 0x1030
    x"F5",x"B6",x"77",x"F1",x"25",x"05",x"C2",x"26", -- 0x1038
    x"B5",x"2C",x"C2",x"21",x"B5",x"C9",x"4C",x"53", -- 0x1040
    x"52",x"45",x"54",x"43",x"41",x"4D",x"4F",x"41", -- 0x1048
    x"44",x"41",x"56",x"45",x"45",x"4E",x"4D",x"52", -- 0x1050
    x"41",x"53",x"59",x"50",x"45",x"4F",x"50",x"59", -- 0x1058
    x"44",x"44",x"52",x"4F",x"44",x"20",x"20",x"28", -- 0x1060
    x"59",x"2F",x"4E",x"29",x"20",x"3F",x"00",x"CD", -- 0x1068
    x"A3",x"B5",x"23",x"EB",x"CD",x"92",x"B5",x"EB", -- 0x1070
    x"36",x"0D",x"21",x"5A",x"F3",x"CD",x"D0",x"BF", -- 0x1078
    x"CD",x"EB",x"BF",x"01",x"00",x"AD",x"C5",x"FE", -- 0x1080
    x"02",x"CA",x"7E",x"B7",x"C1",x"2A",x"4A",x"F3", -- 0x1088
    x"11",x"5A",x"F3",x"EB",x"CD",x"95",x"B5",x"CA", -- 0x1090
    x"1E",x"B4",x"3E",x"20",x"12",x"13",x"05",x"C3", -- 0x1098
    x"87",x"B5",x"2A",x"4A",x"F3",x"06",x"08",x"7E", -- 0x10A0
    x"FE",x"21",x"D8",x"12",x"13",x"23",x"05",x"C2", -- 0x10A8
    x"97",x"B5",x"C9",x"16",x"1E",x"CD",x"23",x"B4", -- 0x10B0
    x"CD",x"61",x"B2",x"11",x"5A",x"F3",x"CD",x"92", -- 0x10B8
    x"B5",x"3E",x"20",x"12",x"0E",x"09",x"CD",x"03", -- 0x10C0
    x"B6",x"36",x"20",x"C9",x"CD",x"76",x"B7",x"C3", -- 0x10C8
    x"00",x"AD",x"E5",x"CD",x"86",x"B4",x"4D",x"44", -- 0x10D0
    x"D1",x"19",x"D8",x"EB",x"CD",x"C1",x"BF",x"CD", -- 0x10D8
    x"6C",x"B6",x"EB",x"C9",x"1B",x"59",x"31",x"3D", -- 0x10E0
    x"44",x"49",x"53",x"4B",x"21",x"00",x"1B",x"59", -- 0x10E8
    x"31",x"3A",x"46",x"49",x"4C",x"45",x"20",x"45", -- 0x10F0
    x"58",x"49",x"53",x"54",x"53",x"21",x"00",x"4C", -- 0x10F8
    x"20",x"00",x"3E",x"20",x"CD",x"F9",x"B5",x"3E", -- 0x1100
    x"08",x"0E",x"0C",x"CD",x"0F",x"F8",x"0D",x"C2", -- 0x1108
    x"FB",x"B5",x"C9",x"21",x"5A",x"F3",x"06",x"FF", -- 0x1110
    x"04",x"7E",x"FE",x"21",x"DA",x"1B",x"B6",x"CD", -- 0x1118
    x"0F",x"F8",x"23",x"C3",x"08",x"B6",x"21",x"5A", -- 0x1120
    x"F3",x"06",x"00",x"11",x"1B",x"B6",x"CD",x"03", -- 0x1128
    x"F8",x"FE",x"0D",x"C8",x"D5",x"FE",x"03",x"CA", -- 0x1130
    x"00",x"AD",x"FE",x"08",x"CA",x"40",x"B6",x"FE", -- 0x1138
    x"7F",x"CA",x"54",x"B6",x"FE",x"20",x"D8",x"CD", -- 0x1140
    x"0F",x"F8",x"77",x"23",x"04",x"78",x"B9",x"C0", -- 0x1148
    x"E5",x"21",x"5D",x"B6",x"CD",x"18",x"F8",x"E1", -- 0x1150
    x"2B",x"05",x"78",x"3C",x"C0",x"04",x"23",x"3E", -- 0x1158
    x"18",x"C3",x"0F",x"F8",x"CD",x"40",x"B6",x"04", -- 0x1160
    x"05",x"C2",x"54",x"B6",x"C9",x"08",x"20",x"08", -- 0x1168
    x"00",x"CD",x"8F",x"B4",x"F5",x"DC",x"00",x"F3", -- 0x1170
    x"F1",x"C3",x"AB",x"B4",x"7C",x"BA",x"C0",x"7D", -- 0x1178
    x"BB",x"C9",x"26",x"16",x"CD",x"3C",x"F8",x"CD", -- 0x1180
    x"89",x"AF",x"21",x"00",x"00",x"E5",x"7E",x"23", -- 0x1188
    x"66",x"6F",x"CD",x"9F",x"B6",x"3E",x"2F",x"CD", -- 0x1190
    x"0F",x"F8",x"E1",x"CD",x"93",x"B6",x"3E",x"48", -- 0x1198
    x"C3",x"0F",x"F8",x"23",x"7E",x"CD",x"15",x"F8", -- 0x11A0
    x"2B",x"7E",x"23",x"23",x"C3",x"15",x"F8",x"AF", -- 0x11A8
    x"4F",x"11",x"F0",x"D8",x"B4",x"F2",x"B3",x"B6", -- 0x11B0
    x"19",x"19",x"19",x"06",x"02",x"CD",x"CD",x"B6", -- 0x11B8
    x"C3",x"B6",x"B6",x"CD",x"CB",x"B6",x"11",x"18", -- 0x11C0
    x"FC",x"CD",x"CB",x"B6",x"11",x"9C",x"FF",x"CD", -- 0x11C8
    x"CB",x"B6",x"1E",x"F6",x"CD",x"CB",x"B6",x"7D", -- 0x11D0
    x"C3",x"DE",x"B6",x"06",x"FF",x"F5",x"04",x"F1", -- 0x11D8
    x"E5",x"19",x"7C",x"A7",x"F2",x"CE",x"B6",x"E1", -- 0x11E0
    x"78",x"B1",x"CA",x"61",x"B2",x"78",x"F6",x"30", -- 0x11E8
    x"4F",x"C3",x"0F",x"F8",x"21",x"4E",x"F3",x"D6", -- 0x11F0
    x"40",x"4F",x"AF",x"3C",x"46",x"23",x"22",x"7B", -- 0x11F8
    x"B6",x"23",x"23",x"0D",x"CA",x"FB",x"B6",x"80", -- 0x1200
    x"C3",x"EB",x"B6",x"21",x"00",x"A0",x"D5",x"EB", -- 0x1208
    x"6F",x"26",x"00",x"29",x"29",x"29",x"29",x"19", -- 0x1210
    x"D1",x"C9",x"CD",x"1B",x"F8",x"FE",x"FF",x"C2", -- 0x1218
    x"18",x"B7",x"32",x"19",x"B7",x"C3",x"0A",x"B7", -- 0x1220
    x"FE",x"00",x"C8",x"32",x"19",x"B7",x"F5",x"C5", -- 0x1228
    x"CD",x"54",x"B7",x"01",x"00",x"30",x"CD",x"66", -- 0x1230
    x"B7",x"05",x"C2",x"26",x"B7",x"C1",x"F1",x"C9", -- 0x1238
    x"CD",x"1B",x"F8",x"3C",x"C2",x"30",x"B7",x"C9", -- 0x1240
    x"0E",x"50",x"C3",x"3F",x"B7",x"0E",x"10",x"CD", -- 0x1248
    x"61",x"B7",x"0C",x"79",x"FE",x"A0",x"C2",x"3F", -- 0x1250
    x"B7",x"CD",x"61",x"B7",x"0D",x"79",x"FE",x"10", -- 0x1258
    x"C2",x"49",x"B7",x"C9",x"F5",x"01",x"28",x"40", -- 0x1260
    x"CD",x"61",x"B7",x"05",x"C2",x"58",x"B7",x"F1", -- 0x1268
    x"C9",x"FB",x"CD",x"66",x"B7",x"F3",x"C5",x"0D", -- 0x1270
    x"C2",x"67",x"B7",x"C1",x"C9",x"1A",x"77",x"23", -- 0x1278
    x"13",x"3C",x"C2",x"6D",x"B7",x"C9",x"16",x"4F", -- 0x1280
    x"21",x"D4",x"B5",x"C3",x"83",x"B7",x"16",x"9F", -- 0x1288
    x"21",x"DE",x"B5",x"E5",x"01",x"1C",x"11",x"21", -- 0x1290
    x"9D",x"CF",x"CD",x"8A",x"B3",x"CD",x"5F",x"B4", -- 0x1298
    x"E1",x"CD",x"18",x"F8",x"CD",x"38",x"B7",x"CD", -- 0x12A0
    x"38",x"B7",x"C3",x"03",x"F8",x"E5",x"01",x"11", -- 0x12A8
    x"2F",x"21",x"E9",x"C0",x"CD",x"8A",x"B3",x"CD", -- 0x12B0
    x"5F",x"B4",x"21",x"08",x"18",x"CD",x"3C",x"F8", -- 0x12B8
    x"CD",x"30",x"B7",x"CD",x"62",x"AF",x"CD",x"0F", -- 0x12C0
    x"F8",x"3E",x"3E",x"CD",x"0F",x"F8",x"E1",x"CD", -- 0x12C8
    x"18",x"F8",x"2A",x"4A",x"F3",x"EB",x"21",x"5A", -- 0x12D0
    x"F3",x"0E",x"08",x"1A",x"77",x"CD",x"0F",x"F8", -- 0x12D8
    x"13",x"23",x"FE",x"20",x"C8",x"0D",x"C2",x"CB", -- 0x12E0
    x"B7",x"36",x"20",x"C3",x"61",x"B2",x"16",x"0F", -- 0x12E8
    x"21",x"EF",x"B5",x"CD",x"9D",x"B7",x"0E",x"0F", -- 0x12F0
    x"CD",x"19",x"B6",x"77",x"21",x"5A",x"F3",x"22", -- 0x12F8
    x"4A",x"F3",x"CD",x"61",x"B6",x"2A",x"4A",x"F3", -- 0x1300
    x"CD",x"D0",x"BF",x"21",x"FD",x"BF",x"E5",x"C3", -- 0x1308
    x"3E",x"F3",x"CD",x"FA",x"BF",x"E5",x"B7",x"F8", -- 0x1310
    x"C3",x"8A",x"AD",x"FF",x"C3",x"18",x"F3",x"C3", -- 0x1318
    x"12",x"F3",x"3E",x"01",x"32",x"00",x"F9",x"72", -- 0x1320
    x"3E",x"00",x"32",x"00",x"F9",x"C9",x"AF",x"47", -- 0x1328
    x"4F",x"C3",x"1D",x"F3",x"3E",x"01",x"01",x"1F", -- 0x1330
    x"1F",x"32",x"00",x"F9",x"21",x"00",x"00",x"39", -- 0x1338
    x"31",x"00",x"F0",x"11",x"00",x"03",x"C5",x"C5", -- 0x1340
    x"C5",x"C5",x"C5",x"C5",x"C5",x"C5",x"1B",x"7A", -- 0x1348
    x"B3",x"C2",x"2A",x"F3",x"F9",x"AF",x"32",x"00", -- 0x1350
    x"F9",x"C9",x"FF",x"16",x"4E",x"CD",x"23",x"B4", -- 0x1358
    x"2A",x"4C",x"F3",x"4C",x"CD",x"3C",x"F8",x"21", -- 0x1360
    x"56",x"B5",x"CD",x"18",x"F8",x"CD",x"03",x"F8", -- 0x1368
    x"FE",x"40",x"DA",x"67",x"B8",x"E6",x"5F",x"FE", -- 0x1370
    x"59",x"C2",x"21",x"B4",x"CD",x"62",x"AF",x"D6", -- 0x1378
    x"41",x"CA",x"21",x"B4",x"C5",x"CD",x"C3",x"B8", -- 0x1380
    x"CD",x"61",x"B6",x"CD",x"1E",x"B4",x"C1",x"0D", -- 0x1388
    x"CD",x"70",x"AF",x"CA",x"84",x"AD",x"3E",x"14", -- 0x1390
    x"91",x"FE",x"01",x"CA",x"BA",x"B8",x"32",x"A3", -- 0x1398
    x"B2",x"79",x"87",x"87",x"81",x"87",x"32",x"99", -- 0x13A0
    x"B2",x"CD",x"8A",x"B2",x"3A",x"79",x"F3",x"4F", -- 0x13A8
    x"3A",x"81",x"F3",x"91",x"FE",x"14",x"DA",x"BA", -- 0x13B0
    x"B8",x"3A",x"7D",x"F3",x"32",x"B6",x"B8",x"3E", -- 0x13B8
    x"12",x"81",x"CD",x"E2",x"B1",x"3E",x"00",x"32", -- 0x13C0
    x"7D",x"F3",x"2A",x"4C",x"F3",x"CD",x"72",x"B6", -- 0x13C8
    x"C3",x"C2",x"B4",x"CD",x"B5",x"B4",x"CD",x"EE", -- 0x13D0
    x"BF",x"C3",x"EB",x"B3",x"AF",x"32",x"97",x"B9", -- 0x13D8
    x"CD",x"62",x"AF",x"32",x"41",x"B9",x"16",x"9F", -- 0x13E0
    x"CD",x"23",x"B4",x"CD",x"E5",x"B1",x"01",x"DE", -- 0x13E8
    x"B8",x"C5",x"CD",x"C8",x"B1",x"26",x"01",x"E5", -- 0x13F0
    x"22",x"4C",x"F3",x"CD",x"19",x"B4",x"3E",x"3C", -- 0x13F8
    x"CD",x"0F",x"F8",x"CD",x"C2",x"B7",x"3E",x"08", -- 0x1400
    x"CD",x"0F",x"F8",x"3E",x"3E",x"CD",x"0F",x"F8", -- 0x1408
    x"CD",x"0A",x"B7",x"E1",x"F5",x"CD",x"16",x"B4", -- 0x1410
    x"F1",x"F5",x"CD",x"EC",x"AD",x"F1",x"FE",x"52", -- 0x1418
    x"C2",x"2E",x"B9",x"32",x"97",x"B9",x"CD",x"A3", -- 0x1420
    x"B5",x"21",x"5A",x"F3",x"3E",x"20",x"BE",x"CA", -- 0x1428
    x"3A",x"B9",x"CD",x"5C",x"AF",x"CD",x"B8",x"B4", -- 0x1430
    x"C2",x"3A",x"B9",x"C3",x"40",x"B9",x"FE",x"0D", -- 0x1438
    x"C0",x"CD",x"5C",x"AF",x"CD",x"B5",x"B4",x"CA", -- 0x1440
    x"40",x"B9",x"CD",x"7E",x"B7",x"C3",x"00",x"AD", -- 0x1448
    x"3E",x"00",x"CD",x"D6",x"BF",x"CD",x"B5",x"B4", -- 0x1450
    x"CD",x"C7",x"BF",x"69",x"60",x"22",x"67",x"B9", -- 0x1458
    x"CD",x"5C",x"AF",x"21",x"10",x"00",x"19",x"22", -- 0x1460
    x"6A",x"B9",x"CD",x"C2",x"B5",x"C5",x"DA",x"BC", -- 0x1468
    x"B5",x"CD",x"A2",x"B4",x"D1",x"D5",x"21",x"00", -- 0x1470
    x"00",x"01",x"00",x"00",x"C5",x"3A",x"41",x"B9", -- 0x1478
    x"CD",x"D6",x"BF",x"CD",x"DC",x"BF",x"23",x"4F", -- 0x1480
    x"CD",x"5C",x"AF",x"EB",x"79",x"CD",x"DF",x"BF", -- 0x1488
    x"23",x"EB",x"C1",x"0B",x"78",x"B1",x"C2",x"6C", -- 0x1490
    x"B9",x"EB",x"3E",x"FF",x"CD",x"DF",x"BF",x"21", -- 0x1498
    x"84",x"AD",x"E3",x"11",x"5A",x"F3",x"3E",x"00", -- 0x14A0
    x"B7",x"C8",x"06",x"08",x"E5",x"3E",x"20",x"CD", -- 0x14A8
    x"DF",x"BF",x"23",x"05",x"C2",x"9D",x"B9",x"E1", -- 0x14B0
    x"06",x"08",x"1A",x"F5",x"CD",x"DF",x"BF",x"F1", -- 0x14B8
    x"23",x"13",x"FE",x"20",x"C8",x"05",x"C2",x"AA", -- 0x14C0
    x"B9",x"C9",x"01",x"30",x"17",x"21",x"7C",x"D0", -- 0x14C8
    x"CD",x"8A",x"B3",x"16",x"0F",x"CD",x"5F",x"B4", -- 0x14D0
    x"21",x"21",x"0D",x"CD",x"3C",x"F8",x"01",x"0C", -- 0x14D8
    x"08",x"16",x"0E",x"CD",x"3B",x"B4",x"21",x"5D", -- 0x14E0
    x"BA",x"CD",x"18",x"F8",x"21",x"1A",x"0F",x"CD", -- 0x14E8
    x"3C",x"F8",x"21",x"62",x"BA",x"CD",x"18",x"F8", -- 0x14F0
    x"CD",x"30",x"B7",x"0E",x"09",x"CD",x"16",x"B6", -- 0x14F8
    x"36",x"20",x"23",x"E5",x"C3",x"FA",x"B9",x"CD", -- 0x1500
    x"55",x"BA",x"21",x"1A",x"10",x"CD",x"3C",x"F8", -- 0x1508
    x"21",x"69",x"BA",x"CD",x"18",x"F8",x"CD",x"F2", -- 0x1510
    x"B5",x"E1",x"E5",x"0E",x"0A",x"CD",x"19",x"B6", -- 0x1518
    x"36",x"0D",x"D1",x"D5",x"CD",x"70",x"BA",x"01", -- 0x1520
    x"F7",x"B9",x"C5",x"C0",x"D8",x"CD",x"6C",x"B6", -- 0x1528
    x"D0",x"C1",x"22",x"50",x"BA",x"01",x"00",x"AD", -- 0x1530
    x"C5",x"E5",x"D5",x"7C",x"2F",x"67",x"7D",x"2F", -- 0x1538
    x"6F",x"19",x"23",x"CD",x"C2",x"B5",x"DA",x"BC", -- 0x1540
    x"B5",x"CD",x"A2",x"B4",x"D1",x"E1",x"CD",x"CA", -- 0x1548
    x"BF",x"21",x"5A",x"F3",x"CD",x"D0",x"BF",x"CD", -- 0x1550
    x"F7",x"BF",x"FE",x"02",x"CA",x"7E",x"B7",x"21", -- 0x1558
    x"00",x"00",x"C3",x"BE",x"BF",x"3E",x"3F",x"CD", -- 0x1560
    x"0F",x"F8",x"C3",x"94",x"B7",x"53",x"41",x"56", -- 0x1568
    x"45",x"00",x"4E",x"41",x"4D",x"45",x"3A",x"20", -- 0x1570
    x"00",x"61",x"44",x"44",x"52",x"3A",x"20",x"00", -- 0x1578
    x"CD",x"7D",x"BA",x"C0",x"D8",x"E5",x"CD",x"7D", -- 0x1580
    x"BA",x"EB",x"E1",x"3F",x"C9",x"21",x"00",x"00", -- 0x1588
    x"C5",x"45",x"4D",x"09",x"1A",x"13",x"FE",x"20", -- 0x1590
    x"CA",x"83",x"BA",x"FE",x"0D",x"CA",x"B5",x"BA", -- 0x1598
    x"FE",x"2C",x"CA",x"B6",x"BA",x"D6",x"30",x"FA", -- 0x15A0
    x"B3",x"BA",x"FE",x"0A",x"FA",x"AB",x"BA",x"FE", -- 0x15A8
    x"11",x"FA",x"B3",x"BA",x"FE",x"17",x"F2",x"B3", -- 0x15B0
    x"BA",x"D6",x"07",x"4F",x"29",x"29",x"29",x"29", -- 0x15B8
    x"D2",x"83",x"BA",x"AF",x"3C",x"37",x"C1",x"C9", -- 0x15C0
    x"CD",x"61",x"B6",x"3E",x"1F",x"CD",x"0F",x"F8", -- 0x15C8
    x"CD",x"B5",x"B4",x"CD",x"CD",x"BF",x"CD",x"DC", -- 0x15D0
    x"BF",x"FE",x"0D",x"C2",x"D6",x"BA",x"CD",x"0F", -- 0x15D8
    x"F8",x"3E",x"0A",x"CD",x"0F",x"F8",x"E6",x"7F", -- 0x15E0
    x"FE",x"7F",x"CA",x"E2",x"BA",x"FE",x"1F",x"D4", -- 0x15E8
    x"0F",x"F8",x"CD",x"1B",x"F8",x"FE",x"03",x"CA", -- 0x15F0
    x"00",x"AD",x"3C",x"C2",x"E2",x"BA",x"23",x"CD", -- 0x15F8
    x"6C",x"B6",x"C2",x"C6",x"BA",x"CD",x"03",x"F8", -- 0x1600
    x"C3",x"00",x"AD",x"00",x"00",x"00",x"00",x"FF", -- 0x1608
    x"53",x"44",x"4F",x"53",x"24",x"20",x"20",x"20", -- 0x1610
    x"00",x"96",x"16",x"08",x"00",x"FF",x"FF",x"FF", -- 0x1618
    x"21",x"16",x"9E",x"01",x"7A",x"A3",x"79",x"95", -- 0x1620
    x"4F",x"78",x"9C",x"47",x"36",x"00",x"23",x"0B", -- 0x1628
    x"79",x"B0",x"C2",x"0C",x"96",x"CD",x"92",x"9B", -- 0x1630
    x"C3",x"00",x"96",x"3E",x"FF",x"32",x"60",x"F7", -- 0x1638
    x"C9",x"3E",x"FF",x"32",x"60",x"F7",x"06",x"0A", -- 0x1640
    x"3E",x"FF",x"32",x"61",x"F7",x"05",x"C2",x"28", -- 0x1648
    x"96",x"3E",x"FE",x"32",x"60",x"F7",x"06",x"10", -- 0x1650
    x"3E",x"40",x"11",x"00",x"00",x"C5",x"CD",x"DB", -- 0x1658
    x"96",x"C1",x"D2",x"51",x"96",x"05",x"C2",x"38", -- 0x1660
    x"96",x"2E",x"00",x"3E",x"FF",x"32",x"60",x"F7", -- 0x1668
    x"C9",x"3E",x"48",x"11",x"AA",x"01",x"CD",x"C2", -- 0x1670
    x"96",x"21",x"A5",x"96",x"DA",x"62",x"96",x"21", -- 0x1678
    x"B3",x"96",x"01",x"78",x"00",x"C5",x"CD",x"7C", -- 0x1680
    x"96",x"C1",x"D2",x"7D",x"96",x"05",x"C2",x"65", -- 0x1688
    x"96",x"0D",x"C2",x"65",x"96",x"3E",x"FF",x"32", -- 0x1690
    x"60",x"F7",x"B7",x"C9",x"E9",x"3E",x"7A",x"11", -- 0x1698
    x"00",x"00",x"CD",x"C2",x"96",x"DA",x"75",x"96", -- 0x16A0
    x"78",x"E6",x"40",x"32",x"BC",x"9D",x"CC",x"9A", -- 0x16A8
    x"96",x"3E",x"FF",x"32",x"60",x"F7",x"3E",x"00", -- 0x16B0
    x"B7",x"C9",x"3E",x"50",x"01",x"00",x"00",x"11", -- 0x16B8
    x"00",x"02",x"C3",x"AC",x"96",x"3E",x"41",x"01", -- 0x16C0
    x"00",x"00",x"50",x"59",x"CD",x"E9",x"96",x"B7", -- 0x16C8
    x"C8",x"37",x"C9",x"3E",x"77",x"CD",x"A7",x"96", -- 0x16D0
    x"3E",x"69",x"01",x"00",x"40",x"51",x"59",x"C3", -- 0x16D8
    x"AC",x"96",x"CD",x"DB",x"96",x"D8",x"F5",x"CD", -- 0x16E0
    x"19",x"97",x"67",x"CD",x"19",x"97",x"6F",x"CD", -- 0x16E8
    x"19",x"97",x"57",x"CD",x"19",x"97",x"5F",x"44", -- 0x16F0
    x"4D",x"F1",x"C9",x"01",x"00",x"00",x"CD",x"E9", -- 0x16F8
    x"96",x"47",x"E6",x"FE",x"78",x"C2",x"B1",x"96", -- 0x1700
    x"C9",x"32",x"61",x"F7",x"F5",x"78",x"00",x"32", -- 0x1708
    x"61",x"F7",x"79",x"00",x"32",x"61",x"F7",x"7A", -- 0x1710
    x"00",x"32",x"61",x"F7",x"7B",x"00",x"32",x"61", -- 0x1718
    x"F7",x"F1",x"FE",x"40",x"06",x"95",x"CA",x"12", -- 0x1720
    x"97",x"FE",x"48",x"06",x"87",x"CA",x"12",x"97", -- 0x1728
    x"06",x"FF",x"78",x"32",x"61",x"F7",x"C3",x"19", -- 0x1730
    x"97",x"01",x"64",x"00",x"3A",x"61",x"F7",x"FE", -- 0x1738
    x"FF",x"C0",x"05",x"C2",x"1C",x"97",x"0D",x"C2", -- 0x1740
    x"1C",x"97",x"C9",x"06",x"00",x"3E",x"FE",x"32", -- 0x1748
    x"60",x"F7",x"3A",x"BC",x"9D",x"B7",x"CC",x"60", -- 0x1750
    x"97",x"3E",x"51",x"CD",x"AC",x"96",x"D2",x"42", -- 0x1758
    x"97",x"C9",x"CD",x"6C",x"97",x"DA",x"41",x"97", -- 0x1760
    x"06",x"00",x"3A",x"61",x"F7",x"00",x"77",x"23", -- 0x1768
    x"3A",x"61",x"F7",x"77",x"23",x"05",x"C2",x"4A", -- 0x1770
    x"97",x"3A",x"61",x"F7",x"3A",x"61",x"F7",x"C9", -- 0x1778
    x"E5",x"EB",x"79",x"29",x"8F",x"47",x"4C",x"55", -- 0x1780
    x"1E",x"00",x"E1",x"C9",x"06",x"FF",x"C5",x"CD", -- 0x1788
    x"19",x"97",x"C1",x"FE",x"FE",x"C8",x"05",x"C2", -- 0x1790
    x"6E",x"97",x"37",x"C9",x"21",x"4E",x"9E",x"7E", -- 0x1798
    x"23",x"FE",x"46",x"C0",x"7E",x"23",x"FE",x"41", -- 0x17A0
    x"C0",x"7E",x"FE",x"54",x"C9",x"AF",x"CD",x"91", -- 0x17A8
    x"97",x"CD",x"94",x"97",x"0A",x"8D",x"12",x"6C", -- 0x17B0
    x"26",x"00",x"03",x"13",x"C9",x"5E",x"23",x"56", -- 0x17B8
    x"23",x"4E",x"23",x"46",x"C9",x"7E",x"83",x"77", -- 0x17C0
    x"23",x"7E",x"8A",x"77",x"23",x"7E",x"89",x"77", -- 0x17C8
    x"23",x"7E",x"88",x"77",x"C9",x"7E",x"83",x"5F", -- 0x17D0
    x"23",x"7E",x"8A",x"57",x"23",x"7E",x"89",x"4F", -- 0x17D8
    x"23",x"7E",x"88",x"47",x"C9",x"7B",x"87",x"5F", -- 0x17E0
    x"7A",x"8F",x"57",x"79",x"8F",x"4F",x"78",x"8F", -- 0x17E8
    x"47",x"C9",x"CD",x"D5",x"97",x"CD",x"D8",x"97", -- 0x17F0
    x"CD",x"DB",x"97",x"0F",x"F5",x"D2",x"E5",x"97", -- 0x17F8
    x"E5",x"CD",x"A5",x"97",x"E1",x"CD",x"C5",x"97", -- 0x1800
    x"F1",x"C9",x"CD",x"EF",x"97",x"C0",x"23",x"34", -- 0x1808
    x"C0",x"23",x"34",x"C9",x"1C",x"C0",x"14",x"C0", -- 0x1810
    x"0C",x"C0",x"04",x"C9",x"13",x"13",x"13",x"23", -- 0x1818
    x"23",x"23",x"CD",x"08",x"98",x"C0",x"1B",x"2B", -- 0x1820
    x"1A",x"96",x"C0",x"1B",x"2B",x"1A",x"96",x"C9", -- 0x1828
    x"7E",x"23",x"B6",x"23",x"B6",x"23",x"B6",x"C9", -- 0x1830
    x"7D",x"91",x"6F",x"7C",x"98",x"67",x"C9",x"01", -- 0x1838
    x"04",x"00",x"79",x"B7",x"CA",x"28",x"98",x"04", -- 0x1840
    x"1A",x"77",x"13",x"23",x"0D",x"C2",x"28",x"98", -- 0x1848
    x"05",x"C2",x"28",x"98",x"C9",x"1A",x"96",x"C0", -- 0x1850
    x"13",x"23",x"0B",x"78",x"B1",x"C2",x"35",x"98", -- 0x1858
    x"C9",x"7E",x"B9",x"C8",x"B7",x"37",x"C8",x"23", -- 0x1860
    x"C3",x"41",x"98",x"1A",x"77",x"B7",x"C8",x"13", -- 0x1868
    x"23",x"C3",x"4B",x"98",x"1A",x"FE",x"61",x"D8", -- 0x1870
    x"FE",x"7B",x"D0",x"E6",x"DF",x"C9",x"0E",x"0B", -- 0x1878
    x"CD",x"54",x"98",x"B7",x"CA",x"8E",x"98",x"FE", -- 0x1880
    x"2E",x"CA",x"7F",x"98",x"FE",x"2A",x"CA",x"98", -- 0x1888
    x"98",x"FE",x"3F",x"CA",x"78",x"98",x"BE",x"C0", -- 0x1890
    x"13",x"23",x"0D",x"C2",x"60",x"98",x"C9",x"79", -- 0x1898
    x"FE",x"0B",x"CA",x"C3",x"98",x"FE",x"04",x"DA", -- 0x18A0
    x"94",x"98",x"C2",x"8E",x"98",x"13",x"3E",x"20", -- 0x18A8
    x"1B",x"C3",x"76",x"98",x"13",x"C3",x"60",x"98", -- 0x18B0
    x"13",x"CD",x"54",x"98",x"B7",x"C8",x"06",x"10", -- 0x18B8
    x"FE",x"2E",x"C2",x"AB",x"98",x"79",x"D6",x"02", -- 0x18C0
    x"47",x"3E",x"20",x"05",x"CA",x"94",x"98",x"BE", -- 0x18C8
    x"CA",x"BA",x"98",x"23",x"0D",x"C2",x"AB",x"98", -- 0x18D0
    x"B7",x"C9",x"1A",x"FE",x"2E",x"CA",x"60",x"98", -- 0x18D8
    x"C3",x"78",x"98",x"1A",x"B7",x"C2",x"CB",x"98", -- 0x18E0
    x"1B",x"3E",x"20",x"BE",x"C0",x"13",x"23",x"0D", -- 0x18E8
    x"C2",x"C3",x"98",x"1A",x"B7",x"C9",x"21",x"2C", -- 0x18F0
    x"A3",x"7E",x"BB",x"C2",x"E8",x"98",x"23",x"7E", -- 0x18F8
    x"BA",x"C2",x"E8",x"98",x"23",x"7E",x"B9",x"C8", -- 0x1900
    x"21",x"2C",x"A3",x"73",x"23",x"72",x"23",x"71", -- 0x1908
    x"21",x"18",x"9E",x"C3",x"2B",x"97",x"CD",x"21", -- 0x1910
    x"96",x"C0",x"11",x"00",x"00",x"4B",x"CD",x"E8", -- 0x1918
    x"98",x"D8",x"CD",x"12",x"99",x"D0",x"2A",x"DE", -- 0x1920
    x"9F",x"EB",x"3A",x"E0",x"9F",x"4F",x"CD",x"E8", -- 0x1928
    x"98",x"D8",x"CD",x"7C",x"97",x"37",x"C0",x"2A", -- 0x1930
    x"26",x"9E",x"01",x"34",x"9E",x"11",x"18",x"A3", -- 0x1938
    x"CD",x"8D",x"97",x"2A",x"2E",x"9E",x"EB",x"2A", -- 0x1940
    x"26",x"9E",x"3A",x"28",x"9E",x"19",x"3D",x"C2", -- 0x1948
    x"2D",x"99",x"01",x"34",x"9E",x"11",x"1C",x"A3", -- 0x1950
    x"CD",x"8D",x"97",x"2A",x"29",x"9E",x"22",x"24", -- 0x1958
    x"A3",x"29",x"8F",x"29",x"8F",x"29",x"8F",x"29", -- 0x1960
    x"8F",x"6C",x"67",x"22",x"26",x"A3",x"01",x"1C", -- 0x1968
    x"A3",x"11",x"20",x"A3",x"CD",x"8D",x"97",x"3A", -- 0x1970
    x"25",x"9E",x"32",x"28",x"A3",x"3E",x"C3",x"32", -- 0x1978
    x"29",x"A3",x"3A",x"52",x"9E",x"FE",x"36",x"CC", -- 0x1980
    x"8F",x"9B",x"21",x"78",x"99",x"22",x"2A",x"A3", -- 0x1988
    x"21",x"5C",x"00",x"22",x"18",x"A2",x"AF",x"C9", -- 0x1990
    x"21",x"36",x"A3",x"CD",x"9D",x"97",x"21",x"18", -- 0x1998
    x"A3",x"CD",x"B5",x"97",x"CD",x"D6",x"98",x"DA", -- 0x19A0
    x"A4",x"99",x"2A",x"35",x"A3",x"26",x"00",x"29", -- 0x19A8
    x"11",x"18",x"9E",x"19",x"5E",x"23",x"56",x"7B", -- 0x19B0
    x"F6",x"07",x"A2",x"3C",x"CA",x"A4",x"99",x"EB", -- 0x19B8
    x"22",x"35",x"A3",x"C9",x"AF",x"6F",x"67",x"22", -- 0x19C0
    x"35",x"A3",x"22",x"37",x"A3",x"C9",x"E5",x"3A", -- 0x19C8
    x"30",x"A3",x"B7",x"C2",x"EF",x"99",x"21",x"35", -- 0x19D0
    x"A3",x"CD",x"10",x"98",x"C2",x"C2",x"99",x"E1", -- 0x19D8
    x"37",x"C9",x"11",x"20",x"A3",x"21",x"31",x"A3", -- 0x19E0
    x"CD",x"1F",x"98",x"01",x"02",x"00",x"21",x"35", -- 0x19E8
    x"A3",x"7E",x"91",x"5F",x"23",x"7E",x"98",x"57", -- 0x19F0
    x"23",x"7E",x"98",x"4F",x"23",x"7E",x"98",x"47", -- 0x19F8
    x"3A",x"28",x"A3",x"21",x"31",x"A3",x"CD",x"D2", -- 0x1A00
    x"97",x"CD",x"78",x"99",x"3A",x"28",x"A3",x"3D", -- 0x1A08
    x"32",x"30",x"A3",x"21",x"31",x"A3",x"5E",x"23", -- 0x1A10
    x"56",x"23",x"4E",x"2B",x"2B",x"CD",x"EA",x"97", -- 0x1A18
    x"E1",x"C9",x"CD",x"AE",x"99",x"C3",x"2B",x"97", -- 0x1A20
    x"3A",x"3D",x"A3",x"B7",x"C2",x"17",x"9A",x"21", -- 0x1A28
    x"18",x"A0",x"CD",x"02",x"9A",x"D8",x"AF",x"6F", -- 0x1A30
    x"26",x"00",x"3C",x"FE",x"10",x"DA",x"21",x"9A", -- 0x1A38
    x"AF",x"32",x"3D",x"A3",x"29",x"29",x"29",x"29", -- 0x1A40
    x"29",x"11",x"18",x"A0",x"19",x"C9",x"D5",x"3A", -- 0x1A48
    x"19",x"A2",x"B7",x"C2",x"48",x"9A",x"CD",x"A4", -- 0x1A50
    x"99",x"11",x"1C",x"A3",x"21",x"31",x"A3",x"CD", -- 0x1A58
    x"1F",x"98",x"3A",x"26",x"A3",x"C3",x"52",x"9A", -- 0x1A60
    x"11",x"3E",x"A3",x"21",x"35",x"A3",x"CD",x"1F", -- 0x1A68
    x"98",x"AF",x"32",x"30",x"A3",x"AF",x"32",x"3D", -- 0x1A70
    x"A3",x"D1",x"D5",x"CD",x"08",x"9A",x"D1",x"D8", -- 0x1A78
    x"E5",x"0E",x"20",x"AF",x"B6",x"23",x"0D",x"C2", -- 0x1A80
    x"64",x"9A",x"E1",x"B7",x"37",x"C8",x"7E",x"FE", -- 0x1A88
    x"E5",x"CA",x"5A",x"9A",x"D5",x"E5",x"CD",x"5E", -- 0x1A90
    x"98",x"E1",x"D1",x"C8",x"C3",x"5A",x"9A",x"11", -- 0x1A98
    x"14",x"00",x"19",x"4E",x"23",x"46",x"11",x"05", -- 0x1AA0
    x"00",x"19",x"5E",x"23",x"56",x"C9",x"1A",x"D6", -- 0x1AA8
    x"5C",x"C2",x"9B",x"9A",x"32",x"19",x"A2",x"13", -- 0x1AB0
    x"1A",x"B7",x"C8",x"D5",x"1A",x"B7",x"CA",x"AA", -- 0x1AB8
    x"9A",x"13",x"D6",x"5C",x"C2",x"9C",x"9A",x"1B", -- 0x1AC0
    x"12",x"13",x"EB",x"D1",x"E5",x"D5",x"CD",x"2E", -- 0x1AC8
    x"9A",x"C1",x"DA",x"C1",x"9A",x"E5",x"11",x"0B", -- 0x1AD0
    x"00",x"19",x"7E",x"E1",x"07",x"07",x"07",x"07", -- 0x1AD8
    x"3F",x"D1",x"D8",x"D5",x"C5",x"CD",x"7F",x"9A", -- 0x1AE0
    x"21",x"3E",x"A3",x"73",x"23",x"72",x"23",x"71", -- 0x1AE8
    x"23",x"70",x"D1",x"21",x"18",x"A2",x"7E",x"23", -- 0x1AF0
    x"47",x"7E",x"B7",x"C2",x"D7",x"9A",x"1A",x"FE", -- 0x1AF8
    x"2E",x"C2",x"FA",x"9A",x"13",x"1A",x"FE",x"2E", -- 0x1B00
    x"C2",x"06",x"9B",x"2B",x"7E",x"36",x"00",x"FE", -- 0x1B08
    x"5C",x"C2",x"EB",x"9A",x"32",x"18",x"A2",x"C3", -- 0x1B10
    x"06",x"9B",x"78",x"FE",x"5C",x"CA",x"03",x"9B", -- 0x1B18
    x"36",x"5C",x"23",x"CD",x"4B",x"98",x"D1",x"1A", -- 0x1B20
    x"B7",x"C2",x"9B",x"9A",x"C9",x"21",x"00",x"00", -- 0x1B28
    x"22",x"3B",x"A3",x"CD",x"2E",x"9A",x"D8",x"CD", -- 0x1B30
    x"7F",x"9A",x"21",x"35",x"A3",x"73",x"23",x"72", -- 0x1B38
    x"23",x"71",x"23",x"70",x"AF",x"32",x"30",x"A3", -- 0x1B40
    x"C9",x"78",x"B1",x"C8",x"E5",x"2A",x"3B",x"A3", -- 0x1B48
    x"7C",x"B5",x"CA",x"50",x"9B",x"CD",x"18",x"98", -- 0x1B50
    x"D2",x"7E",x"9B",x"D1",x"C5",x"2A",x"3B",x"A3", -- 0x1B58
    x"44",x"4D",x"E1",x"CD",x"18",x"98",x"E5",x"2A", -- 0x1B60
    x"39",x"A3",x"EB",x"CD",x"22",x"98",x"C1",x"E5", -- 0x1B68
    x"78",x"FE",x"02",x"D2",x"6C",x"9B",x"C5",x"21", -- 0x1B70
    x"00",x"02",x"22",x"3B",x"A3",x"21",x"18",x"A0", -- 0x1B78
    x"22",x"39",x"A3",x"CD",x"02",x"9A",x"C1",x"E1", -- 0x1B80
    x"D2",x"29",x"9B",x"C9",x"21",x"00",x"00",x"22", -- 0x1B88
    x"3B",x"A3",x"E1",x"C5",x"CD",x"02",x"9A",x"C1", -- 0x1B90
    x"D8",x"05",x"05",x"C3",x"29",x"9B",x"22",x"3B", -- 0x1B98
    x"A3",x"2A",x"39",x"A3",x"EB",x"E1",x"CD",x"22", -- 0x1BA0
    x"98",x"EB",x"22",x"39",x"A3",x"EB",x"C9",x"F5", -- 0x1BA8
    x"F1",x"C9",x"3E",x"1F",x"CD",x"0F",x"F8",x"21", -- 0x1BB0
    x"C5",x"9D",x"CD",x"18",x"F8",x"CD",x"F6",x"98", -- 0x1BB8
    x"CD",x"1B",x"96",x"0E",x"38",x"21",x"42",x"A3", -- 0x1BC0
    x"36",x"00",x"23",x"0D",x"C2",x"A8",x"9B",x"21", -- 0x1BC8
    x"DC",x"9D",x"CD",x"18",x"F8",x"21",x"18",x"A2", -- 0x1BD0
    x"CD",x"18",x"F8",x"0E",x"3E",x"CD",x"09",x"F8", -- 0x1BD8
    x"CD",x"A6",x"9C",x"21",x"A3",x"9B",x"E5",x"21", -- 0x1BE0
    x"F2",x"9D",x"7E",x"B7",x"CA",x"F7",x"9C",x"11", -- 0x1BE8
    x"42",x"A3",x"7E",x"B7",x"CA",x"E1",x"9B",x"1A", -- 0x1BF0
    x"BE",x"C2",x"EB",x"9B",x"13",x"23",x"C3",x"D2", -- 0x1BF8
    x"9B",x"1A",x"B7",x"CA",x"F6",x"9B",x"FE",x"20", -- 0x1C00
    x"CA",x"F6",x"9B",x"7E",x"23",x"B7",x"C2",x"EB", -- 0x1C08
    x"9B",x"23",x"23",x"C3",x"CA",x"9B",x"23",x"5E", -- 0x1C10
    x"23",x"56",x"CD",x"F0",x"9C",x"EB",x"E9",x"4E", -- 0x1C18
    x"23",x"CD",x"09",x"F8",x"05",x"C2",x"FF",x"9B", -- 0x1C20
    x"C9",x"11",x"44",x"A3",x"13",x"1A",x"FE",x"20", -- 0x1C28
    x"CA",x"0C",x"9C",x"B7",x"C2",x"1A",x"9C",x"11", -- 0x1C30
    x"EC",x"9D",x"CD",x"2E",x"9A",x"DA",x"72",x"9C", -- 0x1C38
    x"E5",x"CD",x"1B",x"F8",x"FE",x"FF",x"C2",x"21", -- 0x1C40
    x"9C",x"01",x"0B",x"00",x"09",x"7E",x"E1",x"E6", -- 0x1C48
    x"08",x"C2",x"67",x"9C",x"06",x"08",x"CD",x"FF", -- 0x1C50
    x"9B",x"0E",x"20",x"CD",x"09",x"F8",x"06",x"03", -- 0x1C58
    x"CD",x"FF",x"9B",x"0E",x"20",x"CD",x"09",x"F8", -- 0x1C60
    x"7E",x"E6",x"10",x"CA",x"57",x"9C",x"21",x"F2", -- 0x1C68
    x"9D",x"CD",x"18",x"F8",x"C3",x"64",x"9C",x"7D", -- 0x1C70
    x"C6",x"12",x"6F",x"7E",x"CD",x"15",x"F8",x"2B", -- 0x1C78
    x"7E",x"CD",x"15",x"F8",x"CD",x"F0",x"9C",x"CD", -- 0x1C80
    x"5A",x"9A",x"D2",x"20",x"9C",x"CD",x"1B",x"96", -- 0x1C88
    x"C9",x"E1",x"CD",x"1B",x"96",x"21",x"E1",x"9D", -- 0x1C90
    x"C3",x"18",x"F8",x"21",x"43",x"A3",x"23",x"7E", -- 0x1C98
    x"FE",x"20",x"CA",x"7E",x"9C",x"B7",x"C2",x"92", -- 0x1CA0
    x"9C",x"CD",x"F0",x"9C",x"21",x"18",x"A2",x"C3", -- 0x1CA8
    x"18",x"F8",x"EB",x"CD",x"8E",x"9A",x"CD",x"1B", -- 0x1CB0
    x"96",x"D0",x"21",x"EE",x"9D",x"C3",x"18",x"F8", -- 0x1CB8
    x"CD",x"1B",x"96",x"C3",x"00",x"F8",x"21",x"42", -- 0x1CC0
    x"A3",x"CD",x"03",x"F8",x"FE",x"08",x"CA",x"C9", -- 0x1CC8
    x"9C",x"FE",x"7F",x"CA",x"C9",x"9C",x"FE",x"18", -- 0x1CD0
    x"CA",x"E2",x"9C",x"36",x"00",x"FE",x"0D",x"C8", -- 0x1CD8
    x"77",x"23",x"4F",x"CD",x"09",x"F8",x"C3",x"A9", -- 0x1CE0
    x"9C",x"7D",x"FE",x"42",x"CA",x"A9",x"9C",x"0E", -- 0x1CE8
    x"08",x"CD",x"09",x"F8",x"0E",x"20",x"CD",x"09", -- 0x1CF0
    x"F8",x"0E",x"08",x"CD",x"09",x"F8",x"2B",x"C3", -- 0x1CF8
    x"A9",x"9C",x"7E",x"B7",x"CA",x"A9",x"9C",x"FE", -- 0x1D00
    x"0D",x"CA",x"A9",x"9C",x"23",x"C3",x"C2",x"9C", -- 0x1D08
    x"21",x"D9",x"9D",x"CD",x"18",x"F8",x"C9",x"CD", -- 0x1D10
    x"F0",x"9C",x"21",x"42",x"A3",x"0E",x"2E",x"CD", -- 0x1D18
    x"41",x"98",x"11",x"06",x"9E",x"CD",x"4B",x"98", -- 0x1D20
    x"11",x"42",x"A3",x"CD",x"0D",x"9B",x"D2",x"28", -- 0x1D28
    x"9D",x"21",x"42",x"A3",x"0E",x"2E",x"CD",x"41", -- 0x1D30
    x"98",x"11",x"0B",x"9E",x"CD",x"4B",x"98",x"11", -- 0x1D38
    x"42",x"A3",x"CD",x"0D",x"9B",x"DA",x"72",x"9C", -- 0x1D40
    x"01",x"10",x"00",x"21",x"42",x"A3",x"CD",x"29", -- 0x1D48
    x"9B",x"21",x"4A",x"A3",x"5E",x"23",x"56",x"23", -- 0x1D50
    x"4E",x"23",x"46",x"C3",x"3E",x"9D",x"03",x"EB", -- 0x1D58
    x"E5",x"C5",x"C5",x"7C",x"CD",x"15",x"F8",x"7D", -- 0x1D60
    x"CD",x"15",x"F8",x"0E",x"2C",x"CD",x"09",x"F8", -- 0x1D68
    x"78",x"CD",x"15",x"F8",x"C1",x"79",x"CD",x"15", -- 0x1D70
    x"F8",x"C1",x"CD",x"29",x"9B",x"C3",x"1B",x"96", -- 0x1D78
    x"11",x"44",x"A3",x"CD",x"0D",x"9B",x"DA",x"72", -- 0x1D80
    x"9C",x"01",x"10",x"00",x"21",x"42",x"A3",x"CD", -- 0x1D88
    x"29",x"9B",x"21",x"4A",x"A3",x"5E",x"23",x"56", -- 0x1D90
    x"23",x"4E",x"23",x"46",x"D5",x"C5",x"7A",x"CD", -- 0x1D98
    x"15",x"F8",x"7B",x"CD",x"15",x"F8",x"3E",x"2C", -- 0x1DA0
    x"CD",x"0F",x"F8",x"78",x"CD",x"15",x"F8",x"79", -- 0x1DA8
    x"CD",x"15",x"F8",x"21",x"00",x"00",x"CD",x"29", -- 0x1DB0
    x"9B",x"CD",x"1B",x"96",x"3E",x"42",x"CD",x"D6", -- 0x1DB8
    x"BF",x"21",x"42",x"A3",x"CD",x"D0",x"BF",x"21", -- 0x1DC0
    x"00",x"00",x"D1",x"1B",x"CD",x"CA",x"BF",x"CD", -- 0x1DC8
    x"F7",x"BF",x"E1",x"CD",x"BE",x"BF",x"21",x"10", -- 0x1DD0
    x"9E",x"C3",x"18",x"F8",x"00",x"46",x"41",x"54", -- 0x1DD8
    x"00",x"31",x"36",x"0A",x"00",x"53",x"44",x"4F", -- 0x1DE0
    x"53",x"0D",x"0A",x"4F",x"52",x"49",x"20",x"45", -- 0x1DE8
    x"44",x"49",x"54",x"49",x"4F",x"4E",x"0D",x"0A", -- 0x1DF0
    x"00",x"0D",x"0A",x"00",x"0D",x"0A",x"41",x"3A", -- 0x1DF8
    x"00",x"4E",x"4F",x"20",x"46",x"49",x"4C",x"45", -- 0x1E00
    x"28",x"53",x"29",x"00",x"2A",x"00",x"0D",x"4E", -- 0x1E08
    x"4F",x"20",x"44",x"49",x"52",x"00",x"09",x"9C", -- 0x1E10
    x"43",x"44",x"00",x"7B",x"9C",x"58",x"00",x"A0", -- 0x1E18
    x"9C",x"4C",x"00",x"60",x"9D",x"00",x"2E",x"4F", -- 0x1E20
    x"52",x"44",x"00",x"2E",x"42",x"52",x"55",x"00", -- 0x1E28
    x"0D",x"0A",x"4F",x"4B",x"0D",x"00",x"FF",x"FF", -- 0x1E30
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E38
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00", -- 0x1E40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1ED0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1ED8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FD8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"  -- 0x1FF8
  );

begin

  p_rom : process(clk)
  begin
    if rising_edge(clk) then
      data <= ROM(to_integer(unsigned(addr)));
    end if;
  end process;

end RTL;
